library IEEE;
use IEEE.std_logic_1164.ALL;

entity shiftregister_9bit_tb is
end shiftregister_9bit_tb;

