configuration sendfsm_synthesised_cfg of sendfsm is
   for synthesised
      -- skipping lhqd1bwp7t because it is not a local entity
      -- skipping ao221d0bwp7t because it is not a local entity
      -- skipping oai21d0bwp7t because it is not a local entity
      -- skipping oai221d0bwp7t because it is not a local entity
      -- skipping oa31d0bwp7t because it is not a local entity
      -- skipping invd8bwp7t because it is not a local entity
      -- skipping lhd1bwp7t because it is not a local entity
      -- skipping oa21d0bwp7t because it is not a local entity
      -- skipping an4d1bwp7t because it is not a local entity
      -- skipping an2d4bwp7t because it is not a local entity
      -- skipping invd1bwp7t because it is not a local entity
      -- skipping an2d1bwp7t because it is not a local entity
      -- skipping or2d0bwp7t because it is not a local entity
      -- skipping invd0bwp7t because it is not a local entity
      -- skipping dfkcnd1bwp7t because it is not a local entity
      -- skipping tielbwp7t because it is not a local entity
   end for;
end sendfsm_synthesised_cfg;
