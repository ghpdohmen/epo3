library IEEE;
use IEEE.std_logic_1164.ALL;

architecture behaviour of vga_main is
begin
end behaviour;

