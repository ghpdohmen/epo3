configuration vgatest_tb_behaviour_cfg3 of vgatest_tb is
   for behaviour
      for all: vgatest use configuration work.vgatest_routed_cfg;
      end for;
   end for;
end vgatest_tb_behaviour_cfg3;
