library IEEE;
use IEEE.std_logic_1164.ALL;

architecture behaviour of submod_rom is
-- define the new type for the 1023 rom 
type rom_array is array (0 to M ) of std_logic_vector (1 downto 0);
-- initial values in the rom
signal rom: rom_array :=( --00 zwart, 01 doorzichtig, 10 geel, 11 wit
        "01","01","01", "01", "01",--1
        "01","01","01", "01", "01",
        "01","01","01", "01", "01",
        "01","01","01", "01", "01",
        "01","01","01", "01", "01",
        "00","00","00", "00", "01",
        "01", "01",
        "01","01","01", "01", "01",--2 
        "01","01","01", "01", "01",     
        "01","01","01", "01", "01",     
        "01","01","01", "01", "01",     
        "01","01","01", "01", "00",   
        "00","11","11", "00", "00",
        "00", "01",
        "01","01","01", "01", "01",--3
        "01","01","01", "01", "01",
        "01","01","01", "01", "01",
        "01","01","01", "01", "01",
        "01","01","01", "00", "00",
        "00","11","00", "00", "11",
        "00", "00",
        "01","01","01", "01", "01",--4
        "01","01","01", "01", "01",
        "01","01","01", "01", "01",
        "01","01","01", "01", "01",
        "01","01","00", "10", "10",
        "00","11","00", "00", "00",
        "11", "00",
        "01","01","01", "01", "01",--5
        "01","01","01", "01", "01",
        "01","01","01", "01", "01",
        "01","01","01", "01", "01",
        "01","00","10", "10", "10",
        "00","00","11", "00", "00",
        "11", "00",
        "01","01","01", "01", "01",--6
        "01","01","01", "01", "01",
        "01","01","01", "01", "01",
        "01","01","01", "01", "01",
        "00","10","10", "10", "00",
        "10","00","00", "11", "11",
        "11", "00",
        "01","01","01", "01", "01",--7
        "01","01","01", "01", "01",
        "01","01","01", "01", "01",
        "01","01","01", "01", "00",
        "10","10","10", "00", "10",
        "10","10","00", "00", "00",
        "00", "00",
        "01","01","01", "01", "01",--8
        "01","01","01", "01", "01",
        "01","01","01", "01", "01",
        "01","01","01", "00", "10",
        "10","10","00", "10", "10",
        "10","00","10", "10", "10",
        "00", "01",
        "01","01", "01", "01", --9
        "01","01","01", "01", "01",
        "01","01","01", "01", "01",
        "01","01","01", "00", "10",
        "10","10","00", "10", "10",
        "10","00","10", "10", "10",
        "00", "01","01",
        "01", "01", "01", --10
        "01","01","01", "01", "01",
        "01","01","01", "01", "01",
        "01","01","01", "00", "10",
        "10","10","00", "10", "10",
        "10","00","10", "10", "10",
        "00", "01","01","01",
        "01", "01", --11
        "01","01","01", "01", "01",
        "01","01","01", "01", "01",
        "01","01","01", "00", "10",
        "10","10","00", "10", "10",
        "10","00","10", "10", "10",
        "00", "01","01","01","01",
        "01", --12
        "01","01","01", "01", "01",
        "01","01","01", "01", "01",
        "01","01","01", "00", "10",
        "10","10","00", "10", "10",
        "10","00","10", "10", "10",
        "00", "01","01","01","01",
        "01",
        "01","01","01", "01", "01",--13
        "01","01","01", "01", "01",
        "01","01","01", "00", "10",
        "10","10","00", "10", "10",
        "10","00","10", "10", "10",
        "00", "01","01","01","01",
        "01","01",
        "01","01", "01", "01",--14
        "01","01","01", "01", "01",
        "01","01","01", "00", "10",
        "10","10","00", "10", "10",
        "10","00","10", "10", "10",
        "00", "01","01","01","01",
        "01","01","01",
        "01", "01", "01",--15
        "01","01","01", "01", "01",
        "01","01","01", "00", "10",
        "10","10","00", "10", "10",
        "10","00","10", "10", "10",
        "00", "01","01","01","01",
        "01","01","01","01",
        "01", "01",--16
        "01","01","01", "01", "01",
        "01","01","01", "00", "10",
        "10","10","00", "10", "10",
        "10","00","10", "10", "10",
        "00", "01","01","01","01",
        "01","01","01","01","01",
        "01",--17
        "01","01","01", "01", "01",
        "01","01","01", "00", "10",
        "10","10","00", "10", "10",
        "10","00","10", "10", "10",
        "00", "01","01","01","01",
        "01","01","01","01","01",
        "01",
        "01","01","01", "01", "01",--18
        "01","01","01", "00", "10",
        "10","10","00", "10", "10",
        "10","00","10", "10", "10",
        "00", "01","01","01","01",
        "01","01","01","01","01",
        "01","01",
        "01","01", "01", "01",--19
        "01","01","01", "00", "10",
        "10","10","00", "10", "10",
        "10","00","10", "10", "10",
        "00", "01","01","01","01",
        "01","01","01","01","01",
        "01","01","01",
        "01", "01", "01",--20
        "01","01","01", "00", "10",
        "10","10","00", "10", "10",
        "10","00","10", "10", "10",
        "00", "01","01","01","01",
        "01","01","01","01","01",
        "01","01","01","01",
        "01", "01",--21
        "01","01","01", "00", "10",
        "10","10","00", "10", "10",
        "10","00","10", "10", "10",
        "00", "01","01","01","01",
        "01","01","01","01","01",
        "01","01","01","01","01",
        "01",--22
        "01","01","01", "00", "10",
        "10","10","00", "10", "10",
        "10","00","10", "10", "10",
        "00", "01","01","01","01",
        "01","01","01","01","01",
        "01","01","01","01","01",
        "01",
        "01","01","01", "00", "10",--23
        "10","10","00", "10", "10",
        "10","00","10", "10", "10",
        "00", "01","01","01","01",
        "01","01","01","01","01",
        "01","01","01","01","01",
        "01","01",
        "01","01", "00", "10",--24
        "10","10","00", "10", "10",
        "10","00","10", "10", "10",
        "00", "01","01","01","01",
        "01","01","01","01","01",
        "01","01","01","01","01",
        "01","01","01",
        "01", "00", "10",--25
        "10","10","00", "10", "10",
        "10","00","10", "10", "10",
        "00", "01","01","01","01",
        "01","01","01","01","01",
        "01","01","01","01","01",
        "01","01","01","01",
        "01", "00",--26
        "10","10","00", "10", "10",
        "10","00","10", "10", "10",
        "00", "01","01","01","01",
        "01","01","01","01","01",
        "01","01","01","01","01",
        "01","01","01","01","01",
        "01",--27
        "00","10","00", "10", "10",
        "10","00","10", "10", "10",
        "00", "01","01","01","01",
        "01","01","01","01","01",
        "01","01","01","01","01",
        "01","01","01","01","01",
        "01",    
        "01","00","00", "10", "10",--28
        "10","00","10", "10", "10",
        "00", "01","01","01","01",
        "01","01","01","01","01",
        "01","01","01","01","01",
        "01","01","01","01","01",
        "01","01",
        "01","00", "00", "00",--29
        "10","00","10", "10", "10",
        "00", "01","01","01","01",
        "01","01","01","01","01",
        "01","01","01","01","01",
        "01","01","01","01","01",
        "01","01","01",
        "01", "00", "00",--30
        "00","00","10", "10", "10",
        "00", "01","01","01","01",
        "01","01","01","01","01",
        "01","01","01","01","01",
        "01","01","01","01","01",
        "01","01","01","01",
        "01","00","00", "00", "00",--31
        "00","00","00", "01", "01",
        "01","01","01", "01", "01",
        "01","01","01", "01", "01",
        "01","01","01", "01", "01",
        "01","01","01", "01", "01",
        "01", "01",
        "01","01","01", "01", "01",--32
        "01","01","01", "01", "01",
        "01","01","01", "01", "01",
        "01","01","01", "01", "01",
        "01","01","01", "01", "01",
        "01","01","01", "01", "01",
        "01", "01"
   );
signal rom_asked : integer range 0 to 1023;

begin


rom_asked <= to_integer(unsigned(rom_e_asked));
 -- Data to be read out 
process(clk)
begin
if (clk='1') then
        rom_colour_out <= rom(rom_asked);
end if;
end process;
end behaviour;

