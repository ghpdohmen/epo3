configuration vgadrive_behaviour_cfg of vgadrive is
   for behaviour
   end for;
end vgadrive_behaviour_cfg;
