configuration edge_debounce_behav_cfg of edge_debounce is
   for behav
   end for;
end edge_debounce_behav_cfg;
