configuration shiftregister_11bit_behav_cfg of shiftregister_11bit is
   for behav
   end for;
end shiftregister_11bit_behav_cfg;
