library IEEE;
use IEEE.std_logic_1164.ALL;

entity edge_detector_tb is
end edge_detector_tb;

