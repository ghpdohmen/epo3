configuration timebase_behav_cfg of timebase is
   for behav
   end for;
end timebase_behav_cfg;
