library IEEE;
use IEEE.std_logic_1164.ALL;

entity mouse is
   port(mouseX        : out std_logic_vector(2 downto 0);
        buttons       : out std_logic_vector(4 downto 0);
        mouseY        : out std_logic_vector(2 downto 0);
        Handshake_out : out std_logic;
        DataSwitch    : out std_logic;
        ClkSwitch     : out std_logic;
        Handshake_in  : in  std_logic;
        Data_in       : in  std_logic;
        Clk15k        : in  std_logic;
        clk           : in  std_logic;
        reset         : in  std_logic;
		  rst				 : out std_logic);
end mouse;

