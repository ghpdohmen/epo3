configuration syncunit_behaviour_cfg of syncunit is
   for behaviour
   end for;
end syncunit_behaviour_cfg;
