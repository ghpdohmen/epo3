configuration mouse_timer_behav_cfg of mouse_timer is
   for behav
   end for;
end mouse_timer_behav_cfg;
