library IEEE;
use IEEE.std_logic_1164.ALL;

entity vgadriver_tb is
end vgadriver_tb;

