configuration main_fsm_synthesised_cfg of main_fsm is
   for synthesised
      -- skipping oai32d1bwp7t because it is not a local entity
      -- skipping aoi211xd0bwp7t because it is not a local entity
      -- skipping oai31d0bwp7t because it is not a local entity
      -- skipping oai221d0bwp7t because it is not a local entity
      -- skipping oa32d1bwp7t because it is not a local entity
      -- skipping aoi31d0bwp7t because it is not a local entity
      -- skipping oai22d0bwp7t because it is not a local entity
      -- skipping aoi21d0bwp7t because it is not a local entity
      -- skipping moai22d0bwp7t because it is not a local entity
      -- skipping ao32d1bwp7t because it is not a local entity
      -- skipping cknd4bwp7t because it is not a local entity
      -- skipping iao21d0bwp7t because it is not a local entity
      -- skipping or3d4bwp7t because it is not a local entity
      -- skipping nd2d4bwp7t because it is not a local entity
      -- skipping an2d1bwp7t because it is not a local entity
      -- skipping lhd1bwp7t because it is not a local entity
      -- skipping oa21d0bwp7t because it is not a local entity
      -- skipping aoi22d0bwp7t because it is not a local entity
      -- skipping maoi22d0bwp7t because it is not a local entity
      -- skipping an2d4bwp7t because it is not a local entity
      -- skipping ind2d1bwp7t because it is not a local entity
      -- skipping nr2xd0bwp7t because it is not a local entity
      -- skipping invd4bwp7t because it is not a local entity
      -- skipping nd2d0bwp7t because it is not a local entity
      -- skipping ioa21d1bwp7t because it is not a local entity
      -- skipping an3d4bwp7t because it is not a local entity
      -- skipping inr2d1bwp7t because it is not a local entity
      -- skipping invd0bwp7t because it is not a local entity
      -- skipping nd2d1bwp7t because it is not a local entity
      -- skipping nr2d0bwp7t because it is not a local entity
      -- skipping invd1bwp7t because it is not a local entity
      -- skipping dfd1bwp7t because it is not a local entity
      -- skipping dfkcnd1bwp7t because it is not a local entity
   end for;
end main_fsm_synthesised_cfg;
