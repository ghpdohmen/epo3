configuration mux_synthesised_cfg of mux is
   for synthesised
      -- skipping nd2d4bwp7t because it is not a local entity
      -- skipping nd2d0bwp7t because it is not a local entity
      -- skipping ind2d0bwp7t because it is not a local entity
   end for;
end mux_synthesised_cfg;
