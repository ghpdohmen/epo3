configuration pixelgen_behaviour_cfg of pixelgen is
   for behaviour
   end for;
end pixelgen_behaviour_cfg;
