library IEEE;
use IEEE.std_logic_1164.ALL;

entity graphic_toplvl_tb is
end graphic_toplvl_tb;

