configuration rom_cursor_behavioral_cfg of rom_cursor is
   for behavioral
   end for;
end rom_cursor_behavioral_cfg;
