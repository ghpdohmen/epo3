configuration flipflop_bufr_behav_cfg of flipflop_bufr is
   for behav
   end for;
end flipflop_bufr_behav_cfg;
