configuration edge_detector_behav_cfg of edge_detector is
   for behav
   end for;
end edge_detector_behav_cfg;
