configuration vga_main_behaviour_cfg of vga_main is
   for behaviour
   end for;
end vga_main_behaviour_cfg;
