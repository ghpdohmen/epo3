configuration pixel_synthesised_cfg of pixel is
   for synthesised
      -- skipping nd3d0bwp7t because it is not a local entity
      -- skipping ind4d0bwp7t because it is not a local entity
      -- skipping nr4d0bwp7t because it is not a local entity
      -- skipping oai221d0bwp7t because it is not a local entity
      -- skipping cknd2d1bwp7t because it is not a local entity
      -- skipping aoi22d0bwp7t because it is not a local entity
      -- skipping oai32d1bwp7t because it is not a local entity
      -- skipping nr3d0bwp7t because it is not a local entity
      -- skipping aoi211xd0bwp7t because it is not a local entity
      -- skipping nd2d1bwp7t because it is not a local entity
      -- skipping oai22d0bwp7t because it is not a local entity
      -- skipping inr2d1bwp7t because it is not a local entity
      -- skipping nr2d0bwp7t because it is not a local entity
      -- skipping inr2d0bwp7t because it is not a local entity
      -- skipping nd4d0bwp7t because it is not a local entity
      -- skipping oai21d0bwp7t because it is not a local entity
      -- skipping moai22d0bwp7t because it is not a local entity
      -- skipping nd2d0bwp7t because it is not a local entity
      -- skipping aoi21d0bwp7t because it is not a local entity
      -- skipping oai211d1bwp7t because it is not a local entity
      -- skipping ao21d0bwp7t because it is not a local entity
      -- skipping ioa21d1bwp7t because it is not a local entity
      -- skipping oa21d0bwp7t because it is not a local entity
      -- skipping maoi22d0bwp7t because it is not a local entity
      -- skipping xnr2d1bwp7t because it is not a local entity
      -- skipping cknd2d0bwp7t because it is not a local entity
      -- skipping invd1bwp7t because it is not a local entity
      -- skipping cknd1bwp7t because it is not a local entity
      -- skipping invd0bwp7t because it is not a local entity
      -- skipping an4d1bwp7t because it is not a local entity
      -- skipping ckxor2d0bwp7t because it is not a local entity
      -- skipping lnqd1bwp7t because it is not a local entity
      -- skipping ind2d1bwp7t because it is not a local entity
      -- skipping dfkcnqd1bwp7t because it is not a local entity
      -- skipping ckxor2d1bwp7t because it is not a local entity
      -- skipping dfqd1bwp7t because it is not a local entity
      -- skipping oa32d1bwp7t because it is not a local entity
      -- skipping nr2d1bwp7t because it is not a local entity
      -- skipping inr2xd0bwp7t because it is not a local entity
      -- skipping dfd1bwp7t because it is not a local entity
      -- skipping nr2xd0bwp7t because it is not a local entity
      -- skipping oai31d0bwp7t because it is not a local entity
      -- skipping aoi31d0bwp7t because it is not a local entity
      -- skipping lhqd1bwp7t because it is not a local entity
      -- skipping an4d0bwp7t because it is not a local entity
      -- skipping an2d1bwp7t because it is not a local entity
      -- skipping an2d4bwp7t because it is not a local entity
      -- skipping invd2bwp7t because it is not a local entity
      -- skipping aoi221d0bwp7t because it is not a local entity
      -- skipping fa1d0bwp7t because it is not a local entity
      -- skipping ao22d0bwp7t because it is not a local entity
      -- skipping ha1d0bwp7t because it is not a local entity
      -- skipping ind2d0bwp7t because it is not a local entity
      -- skipping inr3d0bwp7t because it is not a local entity
      -- skipping or2d0bwp7t because it is not a local entity
      -- skipping ckan2d1bwp7t because it is not a local entity
      -- skipping lhcnqd1bwp7t because it is not a local entity
      -- skipping lhcnqd2bwp7t because it is not a local entity
      -- skipping nd2d8bwp7t because it is not a local entity
      -- skipping nd2d5bwp7t because it is not a local entity
      -- skipping nd2d6bwp7t because it is not a local entity
      -- skipping nr2xd4bwp7t because it is not a local entity
      -- skipping nr2xd3bwp7t because it is not a local entity
      -- skipping nd2d1p5bwp7t because it is not a local entity
      -- skipping nd4d4bwp7t because it is not a local entity
      -- skipping nr2xd2bwp7t because it is not a local entity
      -- skipping aoi21d2bwp7t because it is not a local entity
      -- skipping nd2d2bwp7t because it is not a local entity
      -- skipping nd2d3bwp7t because it is not a local entity
      -- skipping aoi21d1bwp7t because it is not a local entity
      -- skipping nr2d1p5bwp7t because it is not a local entity
      -- skipping nr2xd1bwp7t because it is not a local entity
      -- skipping oai21d2bwp7t because it is not a local entity
      -- skipping an2d0bwp7t because it is not a local entity
      -- skipping or2d1bwp7t because it is not a local entity
      -- skipping cknd2d2bwp7t because it is not a local entity
      -- skipping maoi222d0bwp7t because it is not a local entity
      -- skipping ioa21d0bwp7t because it is not a local entity
      -- skipping ao21d1bwp7t because it is not a local entity
      -- skipping lnd1bwp7t because it is not a local entity
      -- skipping nd2d4bwp7t because it is not a local entity
      -- skipping aoi22d2bwp7t because it is not a local entity
      -- skipping ioa21d2bwp7t because it is not a local entity
      -- skipping or2d4bwp7t because it is not a local entity
      -- skipping ind3d1bwp7t because it is not a local entity
      -- skipping iao21d0bwp7t because it is not a local entity
      -- skipping oa31d1bwp7t because it is not a local entity
      -- skipping oa22d0bwp7t because it is not a local entity
      -- skipping ao211d0bwp7t because it is not a local entity
      -- skipping or4d1bwp7t because it is not a local entity
      -- skipping oai31d1bwp7t because it is not a local entity
      -- skipping ao222d0bwp7t because it is not a local entity
      -- skipping aoi32d1bwp7t because it is not a local entity
      -- skipping dfxqd1bwp7t because it is not a local entity
      -- skipping edfkcnqd1bwp7t because it is not a local entity
      -- skipping buffd1bwp7t because it is not a local entity
      -- skipping oai222d0bwp7t because it is not a local entity
      -- skipping maoi222d1bwp7t because it is not a local entity
      -- skipping inr4d0bwp7t because it is not a local entity
      -- skipping dfkcnd1bwp7t because it is not a local entity
      -- skipping edfkcnd1bwp7t because it is not a local entity
      -- skipping oai211d0bwp7t because it is not a local entity
      -- skipping or3d0bwp7t because it is not a local entity
      -- skipping ind3d0bwp7t because it is not a local entity
      -- skipping or3d4bwp7t because it is not a local entity
      -- skipping iinr4d0bwp7t because it is not a local entity
      -- skipping an3d1bwp7t because it is not a local entity
      -- skipping mux2nd0bwp7t because it is not a local entity
      -- skipping mux2d1bwp7t because it is not a local entity
      -- skipping tiehbwp7t because it is not a local entity
   end for;
end pixel_synthesised_cfg;
