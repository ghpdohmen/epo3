configuration mux_behav_cfg of mux is
   for behav
   end for;
end mux_behav_cfg;
