configuration main_fsm_behav_cfg of main_fsm is
   for behav
   end for;
end main_fsm_behav_cfg;
