library IEEE;
use IEEE.std_logic_1164.ALL;

entity shiftregister_11bit_tb is
end shiftregister_11bit_tb;

