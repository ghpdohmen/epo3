configuration vgatest_synthesised_cfg of vgatest is
   for synthesised
      -- skipping or4d4bwp7t because it is not a local entity
      -- skipping or3d4bwp7t because it is not a local entity
      -- skipping ckan2d4bwp7t because it is not a local entity
      -- skipping oai31d0bwp7t because it is not a local entity
      -- skipping nr4d0bwp7t because it is not a local entity
      -- skipping ind3d0bwp7t because it is not a local entity
      -- skipping ind4d0bwp7t because it is not a local entity
      -- skipping aoi31d0bwp7t because it is not a local entity
      -- skipping iao21d0bwp7t because it is not a local entity
      -- skipping cknd1bwp7t because it is not a local entity
      -- skipping or2d0bwp7t because it is not a local entity
      -- skipping nd2d0bwp7t because it is not a local entity
      -- skipping mux2nd0bwp7t because it is not a local entity
      -- skipping nd4d0bwp7t because it is not a local entity
      -- skipping invd0bwp7t because it is not a local entity
      -- skipping lnqd1bwp7t because it is not a local entity
      -- skipping lnd1bwp7t because it is not a local entity
      -- skipping buffd12bwp7t because it is not a local entity
      -- skipping dfcnqd1bwp7t because it is not a local entity
      -- skipping nr2xd0bwp7t because it is not a local entity
      -- skipping maoi22d0bwp7t because it is not a local entity
      -- skipping moai22d0bwp7t because it is not a local entity
      -- skipping ind2d1bwp7t because it is not a local entity
      -- skipping ioa21d1bwp7t because it is not a local entity
      -- skipping nd2d1bwp7t because it is not a local entity
      -- skipping inr2xd0bwp7t because it is not a local entity
      -- skipping ind3d1bwp7t because it is not a local entity
      -- skipping nd3d0bwp7t because it is not a local entity
      -- skipping inr3d0bwp7t because it is not a local entity
      -- skipping iind4d0bwp7t because it is not a local entity
      -- skipping xnr2d1bwp7t because it is not a local entity
      -- skipping dfcnd1bwp7t because it is not a local entity
      -- skipping ckxor2d1bwp7t because it is not a local entity
      -- skipping tielbwp7t because it is not a local entity
   end for;
end vgatest_synthesised_cfg;
