library IEEE;
use IEEE.std_logic_1164.ALL;

entity timebase_tb is
end timebase_tb;

