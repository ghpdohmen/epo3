configuration edge_detector_synthesised_cfg of edge_detector is
   for synthesised
      -- skipping an2d4bwp7t because it is not a local entity
      -- skipping dfd1bwp7t because it is not a local entity
      -- skipping dfqd1bwp7t because it is not a local entity
   end for;
end edge_detector_synthesised_cfg;
