configuration submod_rom_behaviour_cfg of submod_rom is
   for behaviour
   end for;
end submod_rom_behaviour_cfg;
