library IEEE;
use IEEE.std_logic_1164.ALL;

entity mouse_tb is
end mouse_tb;

