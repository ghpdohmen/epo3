library IEEE;
use IEEE.std_logic_1164.ALL;

entity vga_main_tb is
end vga_main_tb;

