configuration shiftregister_9bit_behav_cfg of shiftregister_9bit is
   for behav
   end for;
end shiftregister_9bit_behav_cfg;
