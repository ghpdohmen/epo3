configuration colour_storage_behavioral_cfg of colour_storage is
   for behavioral
   end for;
end colour_storage_behavioral_cfg;
