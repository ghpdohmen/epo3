configuration shiftregister_11bit_synthesised_cfg of shiftregister_11bit is
   for synthesised
      -- skipping edfkcnqd1bwp7t because it is not a local entity
      -- skipping invd1bwp7t because it is not a local entity
      -- skipping invd4bwp7t because it is not a local entity
      -- skipping buffd4bwp7t because it is not a local entity
      -- skipping edfkcnd0bwp7t because it is not a local entity
   end for;
end shiftregister_11bit_synthesised_cfg;
