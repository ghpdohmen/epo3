configuration edge_det_fall_behav_cfg of edge_det_fall is
   for behav
   end for;
end edge_det_fall_behav_cfg;
