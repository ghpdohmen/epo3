configuration vgatest_tb_behaviour_cfg2 of vgatest_tb is
   for behaviour
      for all: vgatest use configuration work.vgatest_synthesised_cfg;
      end for;
   end for;
end vgatest_tb_behaviour_cfg2;
