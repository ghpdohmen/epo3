configuration flipflop_synthesised_cfg of flipflop is
   for synthesised
      -- skipping edfqd0bwp7t because it is not a local entity
      -- skipping buffd4bwp7t because it is not a local entity
   end for;
end flipflop_synthesised_cfg;
