
library ieee;
use ieee.std_logic_1164.all;
--library tcb018gbwp7t;
--use tcb018gbwp7t.all;

architecture routed of pixel is

  component BUFFD1BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL01BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKBD1BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL015BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKBD0BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component BUFFD0BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKBD8BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component BUFFD1P5BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKBD2BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component BUFFD3BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL02BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL0BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL1BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL2BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL3BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKBD10BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKBD6BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKBD12BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component BUFFD4BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL4BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component INVD1BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component IND2D2BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component ND2D2BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component ND2D3BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component IOA21D2BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component AOI21D2BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component CKND2BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component ND2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component CKND2D4BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component CKND2D2BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component INVD8BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component AN2D4BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component ND2D2P5BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component CKND2D3BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component ND2D4BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component INVD2BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component NR2XD1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component ND2D6BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component CKND1BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component INVD3BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component INVD4BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component BUFFD5BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component BUFFD2BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKND4BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component CKND0BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component CKBD4BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKND3BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component CKND8BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component CKBD3BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component IND2D4BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component ND2D5BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component INVD6BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component CKND10BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component ND2D1P5BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component ND4D4BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component INVD1P5BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component ND3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component IND4D0BWP7T
    port(A1, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component NR4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component OAI221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; ZN : out std_logic);
  end component;

  component CKND2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component AOI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI32D1BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component NR3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component AOI211XD0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component OAI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component INR2D1BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component NR2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component INR2D0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component ND4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component OAI21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component MOAI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component ND2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component AOI21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component OAI211D1BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component AO21D0BWP7T
    port(A1, A2, B : in std_logic; Z : out std_logic);
  end component;

  component IOA21D1BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component OA21D0BWP7T
    port(A1, A2, B : in std_logic; Z : out std_logic);
  end component;

  component MAOI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component XNR2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component CKND2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component INVD0BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component AN4D1BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component CKXOR2D0BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component LNQD1BWP7T
    port(D, EN : in std_logic; Q : out std_logic);
  end component;

  component IND2D1BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component DFKCNQD1BWP7T
    port(CN, CP, D : in std_logic; Q : out std_logic);
  end component;

  component CKXOR2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component DFQD1BWP7T
    port(CP, D : in std_logic; Q : out std_logic);
  end component;

  component OA32D1BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component NR2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component INR2XD0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component DFD1BWP7T
    port(CP, D : in std_logic; Q, QN : out std_logic);
  end component;

  component NR2XD0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI31D0BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component AOI31D0BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component LHQD1BWP7T
    port(D, E : in std_logic; Q : out std_logic);
  end component;

  component AN4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component AN2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component INR2D2BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component AN2D2BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component AOI221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; ZN : out std_logic);
  end component;

  component FA1D0BWP7T
    port(A, B, CI : in std_logic; CO, S : out std_logic);
  end component;

  component AO22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component INR2XD2BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component CKAN2D2BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component NR2D2P5BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component HA1D0BWP7T
    port(A, B : in std_logic; CO, S : out std_logic);
  end component;

  component IND2D0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component INR3D0BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OR2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component CKAN2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component LNQD2BWP7T
    port(D, EN : in std_logic; Q : out std_logic);
  end component;

  component LHCNQD2BWP7T
    port(CDN, D, E : in std_logic; Q : out std_logic);
  end component;

  component LHCNQD1BWP7T
    port(CDN, D, E : in std_logic; Q : out std_logic);
  end component;

  component ND2D8BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component NR2XD8BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component NR2XD2BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component NR2D4BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component NR2XD3BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component NR2D2BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component NR2D3BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI21D2BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component AN2XD1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component MAOI222D0BWP7T
    port(A, B, C : in std_logic; ZN : out std_logic);
  end component;

  component INVD5BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component NR2D1P5BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component OR2D2BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component CKAN2D8BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component NR2D5BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component IOA21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component INR2D4BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component LND1BWP7T
    port(D, EN : in std_logic; Q, QN : out std_logic);
  end component;

  component LND2BWP7T
    port(D, EN : in std_logic; Q, QN : out std_logic);
  end component;

  component AOI22D2BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component IND3D1BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component IAO21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component OA31D1BWP7T
    port(A1, A2, A3, B : in std_logic; Z : out std_logic);
  end component;

  component OA22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component AO211D0BWP7T
    port(A1, A2, B, C : in std_logic; Z : out std_logic);
  end component;

  component AN2D0BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component OR4D1BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component OAI31D1BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component AO222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; Z : out std_logic);
  end component;

  component AOI32D1BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component DFXQD1BWP7T
    port(CP, DA, DB, SA : in std_logic; Q : out std_logic);
  end component;

  component EDFKCNQD1BWP7T
    port(CN, CP, D, E : in std_logic; Q : out std_logic);
  end component;

  component OAI222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; ZN : out std_logic);
  end component;

  component MAOI222D1BWP7T
    port(A, B, C : in std_logic; ZN : out std_logic);
  end component;

  component INR4D0BWP7T
    port(A1, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component DFKCND1BWP7T
    port(CN, CP, D : in std_logic; Q, QN : out std_logic);
  end component;

  component EDFKCND1BWP7T
    port(CN, CP, D, E : in std_logic; Q, QN : out std_logic);
  end component;

  component OAI211D0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component OR3D0BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component IND3D0BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OR3XD1BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component IINR4D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AN3D1BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component MUX2ND0BWP7T
    port(I0, I1, S : in std_logic; ZN : out std_logic);
  end component;

  component MUX2D1BWP7T
    port(I0, I1, S : in std_logic; Z : out std_logic);
  end component;

  component TIEHBWP7T
    port(Z : out std_logic);
  end component;

  signal FE_PHN530_sig_logic_y_2, FE_PHN529_sig_logic_y_1, FE_PHN528_sig_logic_y_3, FE_PHN527_sig_logic_x_3, FE_PHN526_gl_ram_n_819 : std_logic;
  signal FE_PHN525_sig_logic_y_2, FE_PHN524_sig_logic_x_3, FE_PHN523_sig_logic_y_3, FE_PHN522_FE_OFN4_gl_ram_n_1111, FE_PHN521_gl_ram_n_1111 : std_logic;
  signal FE_PHN520_gl_ram_n_1111, FE_PHN519_gl_ram_n_819, FE_PHN518_sig_logic_x_3, FE_PHN517_sig_logic_y_1, FE_PHN516_sig_logic_y_3 : std_logic;
  signal FE_PHN515_gl_ram_n_1111, FE_PHN514_sig_logic_x_2, FE_PHN513_sig_logic_x_0, FE_PHN512_sig_logic_x_1, FE_PHN511_ml_ms_tb_n_5 : std_logic;
  signal FE_PHN510_gl_ram_n_1111, FE_PHN509_ml_ms_tb_n_5, FE_PHN508_ml_ms_cnt_n_7, FE_PHN507_ml_ms_cnt_n_9, FE_PHN506_sig_logic_x_1 : std_logic;
  signal FE_PHN505_sig_logic_x_0, FE_PHN504_ml_ms_count15k_1, FE_PHN503_ml_ms_count25M_3, FE_PHN502_ml_ms_cnt_count_1, FE_PHN501_clk15k_in : std_logic;
  signal FE_PHN500_ml_ms_cntD_n_22, FE_PHN499_ml_ms_cntD_n_12, FE_PHN498_ml_ms_cntD_n_13, FE_PHN497_ml_il_x1_input_register_3, FE_PHN496_ml_ms_cnt_n_17 : std_logic;
  signal FE_PHN495_ml_ms_cnt_n_15, FE_PHN494_ml_ms_cnt_n_21, FE_PHN493_ml_ms_cnt_n_22, FE_PHN492_ml_ms_cnt_n_19, FE_PHN491_ml_ms_cntD_n_9 : std_logic;
  signal FE_PHN490_ml_ms_cntD_n_11, FE_PHN489_ml_ms_cntD_n_10, FE_PHN488_ml_ms_ed_n_8, FE_PHN487_gl_ram_n_1111, FE_PHN486_ml_ms_btnflipfloprst : std_logic;
  signal FE_PHN485_ml_il_y1_n_47, FE_PHN484_ml_il_x1_n_47, FE_PHN483_ml_il_y1_input_register_3, FE_PHN482_ml_il_y1_n_48, FE_PHN481_ml_il_x1_n_48 : std_logic;
  signal FE_PHN480_ml_ms_n_58, FE_PHN479_ml_il_y1_n_49, FE_PHN478_ml_ms_mfsm_n_46, FE_PHN477_ml_ms_mfsm_n_45, FE_PHN476_ml_ms_mfsm_n_43 : std_logic;
  signal FE_PHN475_ml_ms_tb_n_6, FE_PHN474_ml_ms_cnt_n_11, FE_PHN473_ml_ms_mfsm_n_29, FE_PHN472_ml_ms_cnt_n_10, FE_PHN471_ml_ms_n_57 : std_logic;
  signal FE_PHN470_ml_ms_n_54, FE_PHN469_ml_ms_n_60, FE_PHN468_gl_vgd_n_64, FE_PHN467_ml_ms_ed_n_2, FE_PHN466_ml_ms_mfsm_n_42 : std_logic;
  signal FE_PHN465_ml_ms_n_25, FE_PHN464_ml_ms_n_34, FE_PHN463_ml_ms_n_31, FE_PHN462_ml_ms_n_24, FE_PHN461_ml_ms_n_26 : std_logic;
  signal FE_PHN460_ml_ms_n_30, FE_PHN459_ml_ms_n_20, FE_PHN458_ml_ms_n_32, FE_PHN457_ml_ms_n_19, FE_PHN456_ml_ms_ed_n_5 : std_logic;
  signal FE_PHN455_sig_logic_x_2, FE_PHN454_ml_ms_mfsm_state_0, FE_PHN453_gl_vgd_horizontal_counter_7, FE_PHN452_ml_ms_mfsm_n_47, FE_PHN451_gl_vgd_horizontal_counter_8 : std_logic;
  signal FE_PHN450_gl_vgd_horizontal_counter_6, FE_PHN449_gl_vgd_horizontal_counter_4, FE_PHN448_gl_vgd_horizontal_counter_2, FE_PHN447_ml_ms_cnt_count_1, FE_PHN446_gl_vgd_horizontal_counter_5 : std_logic;
  signal FE_PHN445_gl_vgd_horizontal_counter_3, FE_PHN444_gl_vgd_horizontal_counter_1, FE_PHN443_ml_ms_mfsm_state_2, FE_PHN442_gl_vgd_vertical_counter_9, FE_PHN441_ml_il_x1_state_0 : std_logic;
  signal FE_PHN440_ml_buttons_mouse_0, FE_PHN439_ml_ms_count25M_5, FE_PHN438_clk15k_in, FE_PHN437_ml_ms_count25M_4, FE_PHN436_ml_ms_count25M_7 : std_logic;
  signal FE_PHN435_gl_vgd_horizontal_counter_0, FE_PHN434_ml_ms_count25M_3, FE_PHN433_gl_vgd_vertical_counter_7, FE_PHN432_gl_vgd_horizontal_counter_9, FE_PHN431_ml_il_x1_state_1 : std_logic;
  signal FE_PHN430_gl_gr_lg_lv_n_11, FE_PHN429_ml_mouseX_2, FE_PHN428_ml_ms_count15k_1, FE_PHN427_ml_ms_count25M_10, FE_PHN426_gl_gr_lg_lv_n_10 : std_logic;
  signal FE_PHN425_ml_ms_mux_select, FE_PHN424_ml_il_y1_state_0, FE_PHN423_gl_vgd_vertical_counter_5, FE_PHN422_ml_ms_count15k_2, FE_PHN421_gl_vgd_vertical_counter_6 : std_logic;
  signal FE_PHN420_ml_buttons_mouse_1, FE_PHN419_gl_vgd_vertical_counter_3, FE_PHN418_gl_vgd_vertical_counter_4, FE_PHN417_ml_ms_count15k_3, FE_PHN416_ml_ms_sfsm_state_0 : std_logic;
  signal FE_PHN415_ml_ms_count25M_6, FE_PHN414_ml_ms_count15k_0, FE_PHN413_gl_sig_scale_h, FE_PHN412_gl_vgd_vertical_counter_0, FE_PHN411_ml_ms_data_sr_11bit_7 : std_logic;
  signal FE_PHN410_gl_vgd_vertical_counter_1, FE_PHN409_gl_vgd_vertical_counter_2, FE_PHN408_ml_ms_count25M_2, FE_PHN407_gl_gr_lg_lh_n_9, FE_PHN406_gl_gr_lg_lh_n_14 : std_logic;
  signal FE_PHN405_gl_gr_lg_lv_n_14, FE_PHN404_data_in, FE_PHN403_gl_gr_lg_lh_n_11, FE_PHN402_ml_il_y1_state_1, FE_PHN401_ml_mouseY_0 : std_logic;
  signal FE_PHN400_gl_gr_lg_lv_n_13, FE_PHN399_ml_ms_cntD_count_1, FE_PHN398_ml_mouseX_0, FE_PHN397_ml_ms_cntD_n_0, FE_PHN396_ml_ms_cnt_n_0 : std_logic;
  signal FE_PHN395_ml_mouseY_1, FE_PHN394_ml_buttons_mouse_2, FE_PHN393_ml_ms_cntD_n_23, FE_PHN392_ml_mouseY_2, FE_PHN391_ml_mouseX_1 : std_logic;
  signal FE_PHN390_ml_ms_sr11_data_out_1_80, FE_PHN389_gl_gr_lg_lh_n_15, FE_PHN388_ml_ms_sr11_data_out_5_84, FE_PHN387_ml_ms_sr11_data_out_0_79, FE_PHN386_ml_ms_data_sr_11bit_2 : std_logic;
  signal FE_PHN385_ml_ms_data_sr_11bit_4, FE_PHN384_ml_ms_count_debounce_11, FE_PHN383_ml_ms_data_sr_11bit_6, FE_PHN382_gl_sig_scale_v, FE_PHN381_ml_buttons_mouse_4 : std_logic;
  signal FE_PHN380_ml_ms_data_sr_11bit_3, FE_PHN379_ml_ms_count_debounce_10, FE_PHN378_ml_ms_cnt_count_0, FE_PHN377_ml_ms_count_debounce_3, FE_PHN376_gl_gr_lg_le_new_count_e_1 : std_logic;
  signal FE_PHN375_ml_ms_count_debounce_4, FE_PHN374_gl_gr_lg_le_new_count_e_6, FE_PHN373_gl_gr_lg_le_new_count_e_8, FE_PHN372_gl_gr_lg_le_new_count_e_9, FE_PHN371_gl_gr_lg_le_new_count_e_7 : std_logic;
  signal FE_PHN370_ml_ms_ed_reg1, FE_PHN369_gl_gr_lg_le_new_count_e_5, FE_PHN368_gl_gr_lg_lv_l_edge_reg1, FE_PHN367_gl_gr_lg_le_new_count_e_0, FE_PHN366_gl_gr_lg_le_new_count_e_3 : std_logic;
  signal FE_PHN365_gl_gr_lg_lh_l_edge_reg1, FE_PHN364_gl_gr_lg_le_new_count_e_4, FE_PHN363_gl_gr_lg_le_new_count_e_2, FE_PHN362_ml_ms_ed_state_1, FE_PHN361_ml_ms_count_debounce_9 : std_logic;
  signal FE_PHN360_ml_ms_count_debounce_8, FE_PHN359_gl_vgd_vertical_counter_8, FE_PHN358_ml_buttons_mouse_3, FE_PHN357_ml_ms_cntD_count_0, FE_PHN356_ml_ms_cntD_count_2 : std_logic;
  signal FE_PSN355_gl_ram_ram_16_2, FE_PSN354_gl_ram_ram_73_2, FE_PSN353_gl_ram_ram_36_2, FE_PSN352_gl_ram_ram_85_2, FE_PSN351_gl_ram_ram_72_2 : std_logic;
  signal FE_PSN350_gl_ram_ram_55_2, FE_PHN349_FE_OFN4_gl_ram_n_1111, FE_PHN348_FE_OFN4_gl_ram_n_1111, FE_PHN347_FE_OFN4_gl_ram_n_1111, FE_PHN346_FE_OFN4_gl_ram_n_1111 : std_logic;
  signal FE_PHN345_FE_OFN4_gl_ram_n_1111, FE_PHN344_FE_OFN4_gl_ram_n_1111, FE_PHN343_FE_OFN4_gl_ram_n_1111, FE_PHN342_FE_OFN4_gl_ram_n_1111, FE_PHN341_FE_OFN4_gl_ram_n_1111 : std_logic;
  signal FE_PHN340_FE_OFN4_gl_ram_n_1111, FE_PHN339_FE_OFN4_gl_ram_n_1111, FE_PHN338_FE_OFN4_gl_ram_n_1111, FE_PHN337_FE_OFN4_gl_ram_n_1111, FE_PHN336_FE_OFN4_gl_ram_n_1111 : std_logic;
  signal FE_PHN335_FE_OFN4_gl_ram_n_1111, FE_PHN334_FE_OFN4_gl_ram_n_1111, FE_PHN333_FE_OFN4_gl_ram_n_1111, FE_PHN332_FE_OFN4_gl_ram_n_1111, FE_PHN331_FE_OFN4_gl_ram_n_1111 : std_logic;
  signal FE_PHN330_FE_OFN4_gl_ram_n_1111, FE_PHN329_FE_OFN4_gl_ram_n_1111, FE_PHN328_FE_OFN4_gl_ram_n_1111, FE_PHN327_FE_OFN4_gl_ram_n_1111, FE_PHN326_FE_OFN4_gl_ram_n_1111 : std_logic;
  signal FE_PHN325_FE_OFN4_gl_ram_n_1111, FE_PHN324_FE_OFN4_gl_ram_n_1111, FE_PHN323_FE_OFN4_gl_ram_n_1111, FE_PHN322_FE_OFN4_gl_ram_n_1111, FE_PHN321_FE_OFN4_gl_ram_n_1111 : std_logic;
  signal FE_PHN320_FE_OFN4_gl_ram_n_1111, FE_PHN319_gl_ram_n_1111, FE_PHN318_gl_ram_n_1111, FE_PHN317_gl_ram_n_1111, FE_PHN316_sig_logic_y_3 : std_logic;
  signal FE_PHN315_sig_logic_x_2, FE_PHN314_sig_logic_x_3, FE_PHN313_gl_ram_n_1111, FE_PHN312_gl_ram_n_1111, FE_PHN311_gl_ram_n_1111 : std_logic;
  signal FE_PHN310_gl_ram_n_1111, FE_PHN309_gl_ram_n_1111, FE_PHN308_gl_ram_n_1111, FE_PHN307_gl_ram_n_1111, FE_PHN306_gl_ram_n_1111 : std_logic;
  signal FE_PHN305_gl_ram_n_1111, FE_PHN304_gl_ram_n_1111, FE_PHN303_gl_ram_n_1111, FE_PHN302_gl_ram_n_1111, FE_PHN301_gl_ram_n_1111 : std_logic;
  signal FE_PHN300_gl_ram_n_1111, FE_PHN299_gl_ram_n_1111, FE_PHN298_gl_ram_n_1111, FE_PHN297_gl_ram_n_1111, FE_PHN296_gl_ram_n_1310 : std_logic;
  signal FE_PHN295_gl_ram_n_1111, FE_PHN294_gl_ram_n_1311, FE_PHN293_sig_logic_x_3, FE_PHN292_gl_ram_n_819, FE_PHN291_gl_ram_n_1310 : std_logic;
  signal FE_PHN290_gl_ram_n_1111, FE_PHN289_gl_ram_n_1111, FE_PHN288_gl_ram_n_1111, FE_PHN287_sig_logic_x_3, FE_PHN286_sig_logic_x_2 : std_logic;
  signal FE_PHN285_gl_ram_n_819, FE_PHN284_gl_ram_n_1310, FE_PHN283_gl_ram_n_1111, FE_PHN282_gl_ram_n_1111, FE_PHN281_gl_ram_n_1111 : std_logic;
  signal FE_PHN280_gl_ram_n_1111, FE_PHN279_gl_ram_n_1111, FE_PHN278_gl_ram_n_1111, FE_PHN277_gl_ram_n_1111, FE_PHN276_gl_ram_n_1111 : std_logic;
  signal FE_OCPN275_gl_ram_ram_9_0, FE_OCPN274_gl_ram_ram_32_1, FE_OCPN273_gl_ram_ram_13_2, FE_OCPN272_gl_ram_ram_43_0, FE_OCPN271_gl_ram_ram_40_2 : std_logic;
  signal FE_OCPN270_gl_ram_ram_24_2, FE_OCPN269_gl_ram_ram_52_0, FE_RN_90_0, FE_RN_89_0, FE_OCPN268_gl_ram_ram_10_0 : std_logic;
  signal FE_OCPN267_gl_ram_ram_63_0, FE_OCPN266_gl_ram_ram_55_0, FE_RN_88_0, FE_RN_87_0, FE_RN_86_0 : std_logic;
  signal FE_RN_85_0, FE_OCPN265_gl_ram_ram_54_0, FE_OCPN264_gl_ram_ram_30_0, FE_OCPN263_gl_ram_ram_4_0, FE_OCPN262_gl_ram_ram_49_0 : std_logic;
  signal FE_OCPN260_gl_ram_ram_2_0, FE_OCPN259_gl_ram_ram_9_0, FE_OCPN257_gl_ram_ram_42_0, FE_OCPN255_gl_ram_ram_15_0, FE_RN_84_0 : std_logic;
  signal FE_RN_83_0, FE_RN_82_0, FE_RN_81_0, FE_RN_80_0, FE_RN_79_0 : std_logic;
  signal FE_RN_78_0, FE_OCPN252_gl_ram_ram_25_2, FE_OCPN250_gl_ram_ram_24_2, FE_OCPN249_gl_ram_ram_48_2, FE_OCPN248_gl_ram_ram_51_2 : std_logic;
  signal FE_OCPN247_gl_ram_ram_41_2, FE_OCPN246_gl_ram_ram_1_2, FE_OCPN245_gl_ram_ram_5_0, FE_OCPN244_gl_ram_ram_29_2, FE_OCPN243_gl_ram_ram_28_0 : std_logic;
  signal FE_OCPN242_gl_ram_ram_55_1, FE_RN_77_0, FE_RN_76_0, FE_RN_75_0, FE_RN_74_0 : std_logic;
  signal FE_RN_73_0, FE_RN_72_0, FE_RN_71_0, FE_RN_70_0, FE_RN_69_0 : std_logic;
  signal FE_OCPN240_gl_ram_ram_53_2, FE_OCPN239_gl_ram_ram_86_2, FE_OCPN238_gl_ram_ram_69_2, FE_OCPN237_gl_ram_ram_75_2, FE_OCPN236_gl_ram_ram_82_2 : std_logic;
  signal FE_OCPN235_gl_ram_ram_73_2, FE_OCPN233_gl_ram_ram_12_1, FE_OCPN231_gl_ram_ram_50_2, FE_OCPN228_gl_ram_ram_72_2, FE_OCPN226_gl_ram_ram_46_2 : std_logic;
  signal FE_OCPN225_gl_ram_ram_80_2, FE_OCPN221_gl_ram_ram_0_2, FE_OCPN219_gl_ram_ram_87_2, FE_OCPN218_gl_ram_ram_71_2, FE_OCPN217_gl_ram_ram_67_2 : std_logic;
  signal FE_OCPN214_gl_ram_ram_18_2, FE_OCPN210_gl_ram_ram_12_2, FE_OCPN208_gl_ram_ram_15_2, FE_OCPN204_gl_ram_ram_79_2, FE_OCPN203_gl_ram_ram_44_2 : std_logic;
  signal FE_OCPN200_gl_ram_ram_47_2, FE_OCPN199_gl_ram_ram_2_2, FE_OCPN198_gl_ram_ram_65_2, FE_OCPN197_gl_ram_ram_8_2, FE_OCPN196_gl_ram_ram_78_2 : std_logic;
  signal FE_OCPN195_gl_ram_ram_23_2, FE_OCPN194_gl_ram_ram_3_2, FE_OCPN193_gl_ram_ram_92_2, FE_OCPN192_gl_ram_ram_77_2, FE_OCPN191_gl_ram_ram_83_2 : std_logic;
  signal FE_OCPN189_gl_ram_ram_52_0, FE_OCPN186_gl_ram_ram_13_0, FE_OCPN184_gl_ram_ram_54_1, FE_RN_68_0, FE_RN_67_0 : std_logic;
  signal FE_RN_66_0, FE_RN_65_0, FE_RN_64_0, FE_RN_63_0, FE_RN_62_0 : std_logic;
  signal FE_OCPN183_gl_ram_ram_5_2, FE_OCPN180_gl_ram_ram_6_2, FE_OCPN179_gl_ram_ram_99_2, FE_RN_61_0, FE_RN_60_0 : std_logic;
  signal FE_RN_59_0, FE_OCPN175_gl_ram_ram_37_0, FE_RN_58_0, FE_OCPN174_gl_ram_ram_0_1, FE_OCPN173_gl_ram_ram_7_2 : std_logic;
  signal FE_RN_57_0, FE_RN_56_0, FE_RN_55_0, FE_RN_54_0, FE_RN_53_0 : std_logic;
  signal FE_RN_52_0, FE_RN_51_0, FE_RN_50_0, FE_RN_49_0, FE_RN_48_0 : std_logic;
  signal FE_RN_47_0, FE_RN_46_0, FE_RN_45_0, FE_RN_44_0, FE_RN_43_0 : std_logic;
  signal FE_RN_42_0, FE_OCPN170_gl_ram_ram_40_0, FE_OCPN169_gl_ram_ram_57_2, FE_OCPN167_gl_ram_n_14, FE_RN_41_0 : std_logic;
  signal FE_RN_40_0, FE_RN_39_0, FE_RN_38_0, FE_RN_37_0, FE_RN_35_0 : std_logic;
  signal FE_OCPN163_gl_ram_ram_21_2, FE_RN_34_0, FE_RN_33_0, FE_RN_32_0, FE_RN_31_0 : std_logic;
  signal FE_RN_30_0, FE_RN_29_0, FE_RN_28_0, FE_RN_27_0, FE_RN_26_0 : std_logic;
  signal FE_OCPN38_gl_ram_ram_98_2, FE_RN_24_0, FE_OCPN37_gl_ram_ram_97_1, FE_OCPN36_gl_ram_ram_98_0, FE_OFN35_V : std_logic;
  signal FE_OFN34_H, FE_OFN33_clk15k_switch, FE_OFN32_logic_1_1_net, FE_OFN31_reset, FE_OFN30_gl_rom_n_18 : std_logic;
  signal FE_OFN29_gl_rom_n_18, FE_OFN28_gl_rom_n_18, FE_OFN27_gl_rom_n_21, FE_OFN26_gl_rom_n_21, FE_OFN25_gl_rom_n_21 : std_logic;
  signal FE_OFN24_gl_rom_n_20, FE_OFN23_gl_rom_n_20, FE_OFN22_gl_rom_n_20, FE_OFN21_gl_rom_n_16, FE_OFN20_gl_rom_n_16 : std_logic;
  signal FE_OFN19_gl_rom_n_16, FE_OFN18_gl_rom_n_16, FE_OFN17_gl_rom_n_16, FE_OFN16_gl_rom_n_22, FE_OFN15_gl_rom_n_22 : std_logic;
  signal FE_OFN14_gl_rom_n_22, FE_OFN13_gl_rom_n_19, FE_OFN12_gl_rom_n_19, FE_OFN11_gl_rom_n_19, FE_OFN10_gl_rom_n_17 : std_logic;
  signal FE_OFN9_gl_rom_n_17, FE_OFN8_gl_rom_n_17, FE_OFN7_gl_rom_n_15, FE_OFN6_gl_rom_n_15, FE_OFN5_gl_rom_n_15 : std_logic;
  signal FE_OFN4_gl_ram_n_1111, CTS_365, CTS_364, CTS_363, CTS_362 : std_logic;
  signal CTS_361, CTS_360, CTS_359, CTS_358, CTS_357 : std_logic;
  signal CTS_356, CTS_355, CTS_354, CTS_353, CTS_352 : std_logic;
  signal CTS_351, CTS_350, CTS_349, CTS_348, CTS_347 : std_logic;
  signal CTS_346, CTS_345, CTS_344, CTS_343, CTS_342 : std_logic;
  signal CTS_341, CTS_340, CTS_339, CTS_338, CTS_337 : std_logic;
  signal CTS_336, CTS_335, CTS_334, CTS_333, CTS_332 : std_logic;
  signal CTS_331, CTS_330, CTS_329, CTS_328, CTS_327 : std_logic;
  signal CTS_326, CTS_325, CTS_324, CTS_323, CTS_322 : std_logic;
  signal CTS_321, CTS_320, CTS_319, CTS_318, CTS_317 : std_logic;
  signal CTS_316, CTS_315, CTS_314, CTS_313, CTS_312 : std_logic;
  signal CTS_311, CTS_310, CTS_309, CTS_308, CTS_307 : std_logic;
  signal CTS_306, CTS_305, CTS_304, CTS_303, CTS_302 : std_logic;
  signal CTS_301, CTS_300, CTS_299, CTS_298, CTS_297 : std_logic;
  signal CTS_296, CTS_295, CTS_294, CTS_293, CTS_292 : std_logic;
  signal CTS_291, CTS_290, CTS_289, CTS_288, CTS_287 : std_logic;
  signal CTS_286, CTS_285, FE_OCPN159_gl_ram_ram_59_2, FE_RN_23_0, FE_RN_21_0 : std_logic;
  signal FE_RN_20_0, FE_RN_19_0, FE_RN_18_0, FE_RN_17_0, FE_RN_16_0 : std_logic;
  signal FE_RN_15_0, FE_RN_14_0, FE_RN_13_0, FE_OCPN151_gl_ram_ram_15_1, FE_OCPN150_gl_ram_ram_23_1 : std_logic;
  signal FE_RN_12_0, FE_RN_11_0, FE_RN_10_0, FE_RN_9_0, FE_RN_8_0 : std_logic;
  signal FE_OCPN148_gl_ram_ram_4_1, FE_OCPN147_gl_ram_ram_6_1, FE_OCPN146_gl_ram_ram_86_1, FE_OCPN145_gl_ram_ram_88_1, FE_OCPN144_gl_ram_ram_87_1 : std_logic;
  signal FE_OCPN143_gl_ram_ram_3_1, FE_OCPN140_gl_ram_ram_89_1, FE_OCPN139_gl_ram_ram_90_1, FE_OCPN136_gl_ram_ram_51_1, FE_OCPN133_gl_ram_ram_76_1 : std_logic;
  signal FE_OCPN130_gl_ram_ram_80_1, FE_OCPN127_gl_ram_ram_81_1, FE_OCPN126_gl_ram_ram_21_1, FE_OCPN125_gl_ram_ram_67_1, FE_OCPN123_gl_ram_ram_85_1 : std_logic;
  signal FE_OCPN119_gl_ram_ram_91_1, FE_OCPN117_gl_ram_ram_92_1, FE_OCPN116_gl_ram_ram_71_1, FE_OCPN111_gl_ram_ram_10_2, FE_OCPN110_gl_ram_ram_77_1 : std_logic;
  signal FE_OCPN108_gl_ram_ram_76_2, FE_OCPN107_gl_ram_ram_78_1, FE_OCPN103_gl_ram_ram_13_2, FE_OCPN102_gl_ram_ram_79_1, FE_RN_7_0 : std_logic;
  signal FE_OCPN89_gl_ram_ram_24_0, FE_OCPN85_gl_ram_ram_14_2, FE_OCPN77_gl_ram_ram_32_2, FE_OCPN74_gl_ram_ram_21_0, FE_OCPN72_gl_ram_ram_8_1 : std_logic;
  signal FE_OCPN71_gl_ram_ram_1_1, FE_OCPN70_gl_ram_ram_73_1, FE_OCPN67_gl_ram_ram_77_0, FE_RN_6_0, FE_OCPN66_gl_ram_ram_29_0 : std_logic;
  signal FE_OCPN65_gl_ram_ram_74_1, FE_OCPN63_gl_ram_ram_31_0, FE_OCPN61_gl_ram_ram_55_2, FE_OCPN56_gl_ram_ram_33_1, FE_OCPN54_gl_ram_ram_48_1 : std_logic;
  signal FE_OCPN46_gl_ram_ram_41_0, FE_OCPN43_gl_ram_ram_56_0, FE_OCPN42_gl_ram_ram_60_0, FE_OCPN38_gl_ram_ram_48_0, FE_OCPN28_gl_ram_ram_10_1 : std_logic;
  signal FE_OCPN14_gl_ram_ram_28_1, FE_OCPN10_gl_ram_ram_25_1, FE_OCPN8_gl_ram_ram_47_1, FE_RN_5_0, FE_OCPN7_gl_ram_ram_40_1 : std_logic;
  signal FE_OCPN6_gl_ram_ram_30_1, FE_OCPN2_gl_ram_ram_41_1, FE_RN_3_0, FE_OCPN3_gl_ram_n_1448, FE_OCPN2_gl_ram_n_1448 : std_logic;
  signal FE_OCPN1_gl_ram_n_1448, FE_OCPN0_gl_ram_n_1448, FE_RN_2_0, FE_RN_1_0, FE_RN_0_0 : std_logic;
  signal FE_DBTN0_reset : std_logic;
  signal gl_sig_y : std_logic_vector(3 downto 0);
  signal gl_sig_ram : std_logic_vector(2 downto 0);
  signal sig_output_color : std_logic_vector(2 downto 0);
  signal gl_sig_x : std_logic_vector(3 downto 0);
  signal gl_sig_rom : std_logic_vector(1 downto 0);
  signal sig_logic_x : std_logic_vector(3 downto 0);
  signal sig_logic_y : std_logic_vector(3 downto 0);
  signal gl_gr_lg_le_new_count_e : std_logic_vector(9 downto 0);
  signal gl_sig_e : std_logic_vector(9 downto 0);
  signal gl_rom_rom_584 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_587 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_840 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_843 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_257 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_261 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1002 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1007 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1001 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1005 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_256 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_259 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1004 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1003 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_948 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_946 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1000 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1006 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_753 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_757 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_985 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_989 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_988 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_990 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_838 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_839 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_374 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_375 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_986 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_987 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_984 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_991 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_836 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_834 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_372 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_370 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_994 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_999 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_996 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_998 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_369 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_373 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_997 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_995 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_368 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_371 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_992 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_993 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_833 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_837 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1010 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1015 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_752 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_755 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1012 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1014 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_342 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_343 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_832 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_835 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1013 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1011 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1008 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1009 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_340 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_338 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_978 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_983 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_980 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_982 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_337 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_341 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_977 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_981 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_979 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_336 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_339 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_976 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_945 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_949 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_969 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_973 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_726 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_727 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_972 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_974 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_350 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_351 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_970 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_971 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_968 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_975 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_348 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_346 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_638 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_639 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_962 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_967 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_345 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_349 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_964 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_966 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_724 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_722 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_965 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_963 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_960 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_961 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_344 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_347 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_953 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_959 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_636 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_634 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_944 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_947 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_954 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_957 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_358 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_359 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_956 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_958 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_633 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_637 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_356 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_354 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_952 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_955 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_632 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_635 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_937 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_941 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_353 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_357 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_940 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_942 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_938 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_943 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_936 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_939 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_951 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_352 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_355 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_721 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_725 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_382 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_383 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_622 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_623 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_950 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_380 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_378 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_720 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_723 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_914 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_919 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_913 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_917 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_377 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_381 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_916 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_915 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_376 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_379 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_912 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_918 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_620 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_618 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_922 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_927 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_924 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_926 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_366 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_367 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_617 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_621 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_925 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_923 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_364 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_362 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_920 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_921 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_929 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_933 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_616 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_619 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_361 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_365 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_932 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_934 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_360 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_363 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_930 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_931 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_928 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_935 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_905 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_909 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_908 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_910 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_334 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_335 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_729 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_733 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_906 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_911 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_904 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_907 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_332 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_330 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_898 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_903 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_630 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_631 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_329 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_333 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_897 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_901 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_628 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_626 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_328 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_331 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_900 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_899 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_896 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_902 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_732 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_734 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_694 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_695 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_326 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_327 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_692 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_690 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_625 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_629 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_689 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_693 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_688 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_691 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_324 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_322 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_321 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_325 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_662 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_663 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_624 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_627 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_660 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_658 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_320 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_323 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_657 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_661 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_656 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_659 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_730 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_731 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_665 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_671 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_666 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_669 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_122 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_127 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_668 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_670 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_664 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_667 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_593 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_597 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_124 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_126 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_674 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_679 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_728 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_735 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_673 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_677 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_596 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_598 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_125 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_123 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_120 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_121 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_676 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_675 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_672 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_678 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_697 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_701 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_594 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_595 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_700 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_702 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_110 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_111 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_108 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_106 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_698 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_699 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_696 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_703 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_681 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_685 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_592 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_599 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_105 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_109 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_684 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_686 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_682 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_683 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_104 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_107 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_680 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_687 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_737 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_743 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_654 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_655 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_652 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_650 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_89 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_93 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_649 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_653 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_92 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_94 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_648 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_651 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_606 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_607 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_604 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_602 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_642 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_647 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_90 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_91 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_644 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_646 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_645 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_643 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_640 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_641 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_562 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_567 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_88 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_95 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_738 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_741 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_102 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_103 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_564 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_566 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_601 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_605 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_565 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_563 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_100 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_98 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_560 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_561 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_97 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_101 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_530 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_535 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_600 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_603 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_532 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_534 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_533 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_531 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_96 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_99 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_528 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_529 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_740 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_742 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_537 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_541 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_736 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_739 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_540 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_542 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_118 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_119 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_614 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_615 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_538 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_539 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_116 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_114 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_536 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_543 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_546 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_551 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_113 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_117 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_548 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_550 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_612 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_610 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_549 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_547 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_544 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_545 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_112 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_115 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_569 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_573 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_609 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_613 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_86 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_87 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_572 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_574 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_84 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_82 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_570 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_575 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_568 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_571 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_558 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_559 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_608 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_611 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_81 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_85 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_556 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_554 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_80 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_83 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_553 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_557 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_552 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_555 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_522 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_527 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_718 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_719 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_524 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_526 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_78 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_79 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_525 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_523 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_590 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_591 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_520 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_521 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_76 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_74 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_514 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_519 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_73 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_77 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_516 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_518 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_72 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_75 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_517 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_515 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_512 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_513 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_588 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_586 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_70 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_71 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_585 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_589 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_506 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_511 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_505 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_509 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_716 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_714 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_68 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_66 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_508 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_507 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_504 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_510 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_65 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_69 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1016 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1019 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_64 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_67 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_490 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_495 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_489 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_493 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_713 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_717 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_492 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_491 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_488 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_494 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_474 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_479 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_582 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_583 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_476 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_478 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_477 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_475 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_472 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_473 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_580 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_578 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_481 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_485 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_484 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_486 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_482 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_483 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_480 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_487 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_497 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_501 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_712 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_715 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_577 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_581 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_500 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_502 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_498 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_499 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_576 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_579 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_496 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_503 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_465 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_469 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_468 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_470 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_466 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_471 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1020 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1022 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_710 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_711 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_464 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_467 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_457 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_461 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_460 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_462 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_458 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_459 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_456 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_463 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_708 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_706 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_450 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_455 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_452 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_454 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_453 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_451 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_448 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_449 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_441 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_445 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_444 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_446 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_442 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_443 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_440 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_447 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_705 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_709 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_430 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_431 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_428 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_426 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_425 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_429 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_424 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_427 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_704 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_707 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_409 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_413 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_412 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_414 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_410 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_411 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_408 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_415 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_417 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_421 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_420 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_422 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_418 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_423 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_416 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_419 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_433 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_437 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_436 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_438 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_434 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_435 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_432 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_439 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_406 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_407 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_404 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_402 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_401 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_405 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_400 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_403 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_398 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_399 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_396 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_394 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_393 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_397 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_392 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_395 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_385 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_389 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_830 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_831 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_388 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_390 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_386 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_391 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_384 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_387 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_828 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_826 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_825 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_829 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_824 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_827 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_814 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_815 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_812 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_810 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_809 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_813 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_808 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_811 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_822 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_823 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_218 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_223 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_820 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_818 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_220 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_222 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_221 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_219 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_216 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_217 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_756 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_758 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_226 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_229 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_228 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_230 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_224 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_227 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_242 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_247 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_244 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_246 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_817 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_821 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_185 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_189 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_245 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_243 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_188 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_190 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_240 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_241 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_210 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_215 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_186 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_187 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_212 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_214 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_213 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_211 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_184 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_191 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_208 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_209 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_816 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_819 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_254 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_255 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_252 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_250 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_174 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_175 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_172 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_170 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_249 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_253 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_248 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_251 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_238 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_239 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_169 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_173 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_236 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_234 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_168 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_171 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_233 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_237 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_232 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_235 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_201 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_205 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_204 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_206 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_178 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_183 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_790 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_791 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_202 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_203 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_200 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_207 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_177 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_181 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_198 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_199 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_180 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_179 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_196 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_194 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_176 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_182 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_193 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_197 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_192 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_195 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_788 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_786 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_306 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_311 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_146 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_151 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_308 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_310 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_309 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_307 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_148 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_150 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_304 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_305 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_274 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_279 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_149 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_147 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_276 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_278 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_144 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_145 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_277 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_275 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_272 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_273 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_282 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_287 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_785 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_789 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_284 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_286 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_158 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_159 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_285 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_283 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_784 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_787 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_156 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_154 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_280 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_281 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_290 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_295 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_292 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_294 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_153 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_157 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_293 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_291 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_152 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_155 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_288 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_289 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_313 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_317 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_161 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_165 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_316 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_318 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_314 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_315 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_164 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_166 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_312 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_319 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_297 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_301 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_162 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_163 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_300 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_302 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_298 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_299 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_160 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_167 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_296 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_303 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_265 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_269 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_137 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_141 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_268 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_270 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_266 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_267 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_798 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_799 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_140 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_142 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_264 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_271 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_258 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_263 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_138 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_139 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_260 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_262 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_136 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_143 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_130 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_135 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_796 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_794 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_129 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_133 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_132 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_131 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_128 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_134 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_793 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_797 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_62 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_63 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_60 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_58 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_57 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_61 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_56 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_59 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_792 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_795 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_46 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_47 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_44 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_42 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_41 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_45 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_40 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_43 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1021 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_806 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_807 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_54 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_55 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_52 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_50 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_49 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_53 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_48 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_51 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_804 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_802 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_17 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_21 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_20 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_22 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_18 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_19 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_16 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_23 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_25 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_29 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_801 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_805 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_30 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_31 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_28 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_26 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_27 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_24 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_33 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_37 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_36 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_38 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_800 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_803 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_34 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_35 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_32 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_39 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_9 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_13 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_14 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_15 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_12 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_10 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_11 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_777 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_781 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_8 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_2 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_7 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_4 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_6 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_780 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_782 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_5 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_3 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_0 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_778 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_779 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_754 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_759 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_225 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_231 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_776 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_783 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_774 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_775 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_772 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_770 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_769 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_773 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_762 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_767 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_764 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_766 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_768 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_771 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_765 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_763 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_760 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_761 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_745 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_749 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_748 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_750 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_746 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_751 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_744 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_747 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_886 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_887 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_884 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_882 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_881 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_885 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_880 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_883 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_854 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_855 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_852 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_850 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_849 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_853 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1017 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_848 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_851 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_857 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_863 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_858 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_861 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_890 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_895 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_892 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_894 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_860 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_862 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_893 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_891 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_888 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_889 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_856 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_859 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_874 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_879 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_876 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_878 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_877 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_875 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_872 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_873 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_870 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_871 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_866 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_868 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_869 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_867 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_864 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_865 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_841 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_845 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_844 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_846 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_842 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_847 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1018 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1023 : std_logic_vector(1 downto 0);
  signal gl_ram_ram_86 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_87 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_98 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_97 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_96 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_99 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_60 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_61 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_62 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_63 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_59 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_56 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_58 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_57 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_52 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_53 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_51 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_48 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_54 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_55 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_36 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_37 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_50 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_49 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_34 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_33 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_44 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_45 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_42 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_41 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_38 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_39 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_46 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_47 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_43 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_40 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_35 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_32 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_84 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_85 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_28 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_29 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_30 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_31 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_94 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_95 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_80 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_81 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_24 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_25 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_27 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_26 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_12 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_13 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_14 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_15 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_11 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_8 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_82 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_83 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_10 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_9 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_20 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_21 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_22 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_23 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_16 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_17 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_18 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_19 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_76 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_77 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_4 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_5 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_2 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_1 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_6 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_7 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_3 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_0 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_92 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_93 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_75 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_72 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_78 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_79 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_91 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_88 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_90 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_89 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_68 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_69 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_67 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_64 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_74 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_73 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_70 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_71 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_66 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_65 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_position : std_logic_vector(6 downto 0);
  signal gl_ram_x_grid : std_logic_vector(6 downto 0);
  signal gl_ram_y_grid : std_logic_vector(6 downto 0);
  signal ml_ms_sfsm_state : std_logic_vector(3 downto 0);
  signal ml_ms_sr_new_new_data : std_logic_vector(8 downto 0);
  signal ml_ms_count25M : std_logic_vector(12 downto 0);
  signal ml_ms_data_sr_11bit : std_logic_vector(10 downto 0);
  signal ml_ms_btns : std_logic_vector(4 downto 0);
  signal ml_ms_mouse_x : std_logic_vector(2 downto 0);
  signal ml_ms_mouse_y : std_logic_vector(2 downto 0);
  signal ml_ms_mfsm_state : std_logic_vector(4 downto 0);
  signal ml_ms_count15k : std_logic_vector(3 downto 0);
  signal ml_buttons_mouse : std_logic_vector(4 downto 0);
  signal ml_mouseX : std_logic_vector(2 downto 0);
  signal ml_mouseY : std_logic_vector(2 downto 0);
  signal ml_il_y1_input_register : std_logic_vector(3 downto 0);
  signal ml_il_y1_cmbsop_sel : std_logic_vector(1 downto 0);
  signal ml_il_y1_state : std_logic_vector(1 downto 0);
  signal ml_ms_cnt_count : std_logic_vector(12 downto 0);
  signal ml_il_color1_state : std_logic_vector(2 downto 0);
  signal ml_il_color1_next_state : std_logic_vector(2 downto 0);
  signal gl_vgd_horizontal : std_logic_vector(9 downto 0);
  signal gl_vgd_vertical : std_logic_vector(9 downto 0);
  signal gl_vgd_horizontal_counter : std_logic_vector(9 downto 0);
  signal gl_vgd_vertical_counter : std_logic_vector(9 downto 0);
  signal ml_il_x1_input_register : std_logic_vector(3 downto 0);
  signal ml_il_x1_cmbsop_sel : std_logic_vector(1 downto 0);
  signal ml_il_x1_state : std_logic_vector(1 downto 0);
  signal ml_ms_ed_state : std_logic_vector(1 downto 0);
  signal ml_ms_count_debounce : std_logic_vector(12 downto 0);
  signal ml_ms_cntD_count : std_logic_vector(12 downto 0);
  signal UNCONNECTED, UNCONNECTED0, UNCONNECTED1, UNCONNECTED2, UNCONNECTED3 : std_logic;
  signal UNCONNECTED4, UNCONNECTED5, UNCONNECTED6, UNCONNECTED7, UNCONNECTED8 : std_logic;
  signal UNCONNECTED9, UNCONNECTED10, UNCONNECTED11, UNCONNECTED12, UNCONNECTED13 : std_logic;
  signal UNCONNECTED14, UNCONNECTED15, UNCONNECTED16, UNCONNECTED17, gl_gr_lg_le_n_0 : std_logic;
  signal gl_gr_lg_le_n_1, gl_gr_lg_le_n_2, gl_gr_lg_le_n_3, gl_gr_lg_le_n_4, gl_gr_lg_le_n_5 : std_logic;
  signal gl_gr_lg_le_n_6, gl_gr_lg_le_n_7, gl_gr_lg_le_n_8, gl_gr_lg_le_n_9, gl_gr_lg_le_n_10 : std_logic;
  signal gl_gr_lg_le_n_11, gl_gr_lg_le_n_12, gl_gr_lg_le_n_13, gl_gr_lg_le_n_14, gl_gr_lg_le_n_15 : std_logic;
  signal gl_gr_lg_le_n_16, gl_gr_lg_le_n_17, gl_gr_lg_le_n_18, gl_gr_lg_le_n_19, gl_gr_lg_le_n_20 : std_logic;
  signal gl_gr_lg_le_n_21, gl_gr_lg_le_n_22, gl_gr_lg_le_n_23, gl_gr_lg_le_n_24, gl_gr_lg_le_n_25 : std_logic;
  signal gl_gr_lg_le_n_26, gl_gr_lg_le_n_27, gl_gr_lg_le_n_28, gl_gr_lg_le_n_29, gl_gr_lg_le_n_31 : std_logic;
  signal gl_gr_lg_le_n_32, gl_gr_lg_lh_l_edge_n_0, gl_gr_lg_lh_l_edge_reg1, gl_gr_lg_lh_l_edge_reg2, gl_gr_lg_lh_n_0 : std_logic;
  signal gl_gr_lg_lh_n_1, gl_gr_lg_lh_n_2, gl_gr_lg_lh_n_3, gl_gr_lg_lh_n_4, gl_gr_lg_lh_n_5 : std_logic;
  signal gl_gr_lg_lh_n_6, gl_gr_lg_lh_n_7, gl_gr_lg_lh_n_8, gl_gr_lg_lh_n_9, gl_gr_lg_lh_n_10 : std_logic;
  signal gl_gr_lg_lh_n_11, gl_gr_lg_lh_n_12, gl_gr_lg_lh_n_13, gl_gr_lg_lh_n_14, gl_gr_lg_lh_n_15 : std_logic;
  signal gl_gr_lg_lh_sig_edges, gl_gr_lg_lv_l_edge_n_0, gl_gr_lg_lv_l_edge_reg1, gl_gr_lg_lv_l_edge_reg2, gl_gr_lg_lv_n_0 : std_logic;
  signal gl_gr_lg_lv_n_1, gl_gr_lg_lv_n_2, gl_gr_lg_lv_n_3, gl_gr_lg_lv_n_4, gl_gr_lg_lv_n_5 : std_logic;
  signal gl_gr_lg_lv_n_6, gl_gr_lg_lv_n_7, gl_gr_lg_lv_n_8, gl_gr_lg_lv_n_9, gl_gr_lg_lv_n_10 : std_logic;
  signal gl_gr_lg_lv_n_11, gl_gr_lg_lv_n_12, gl_gr_lg_lv_n_13, gl_gr_lg_lv_n_14, gl_gr_lg_lv_sig_edges : std_logic;
  signal gl_gr_lg_sig_countdown_1_145, gl_gr_lg_sig_countdown_2_144, gl_gr_lg_sig_countdown_3_143, gl_gr_lg_sig_countdown_4_142, gl_gr_lg_sig_countdown_5_141 : std_logic;
  signal gl_gr_lg_sig_countdown_6_140, gl_gr_lg_sig_countdown_7_139, gl_n_0, gl_n_1, gl_n_2 : std_logic;
  signal gl_n_3, gl_n_4, gl_n_5, gl_n_6, gl_n_7 : std_logic;
  signal gl_n_8, gl_n_9, gl_n_10, gl_n_11, gl_n_12 : std_logic;
  signal gl_n_14, gl_n_15, gl_n_16, gl_n_18, gl_n_19 : std_logic;
  signal gl_n_20, gl_n_21, gl_n_22, gl_n_23, gl_n_24 : std_logic;
  signal gl_n_25, gl_n_26, gl_n_27, gl_n_28, gl_n_29 : std_logic;
  signal gl_n_30, gl_n_31, gl_n_32, gl_n_33, gl_n_34 : std_logic;
  signal gl_n_35, gl_n_36, gl_n_37, gl_n_38, gl_n_39 : std_logic;
  signal gl_n_40, gl_n_41, gl_n_42, gl_n_43, gl_n_44 : std_logic;
  signal gl_n_45, gl_ram_n_2, gl_ram_n_3, gl_ram_n_4, gl_ram_n_5 : std_logic;
  signal gl_ram_n_6, gl_ram_n_7, gl_ram_n_8, gl_ram_n_9, gl_ram_n_11 : std_logic;
  signal gl_ram_n_14, gl_ram_n_15, gl_ram_n_16, gl_ram_n_17, gl_ram_n_18 : std_logic;
  signal gl_ram_n_19, gl_ram_n_20, gl_ram_n_21, gl_ram_n_22, gl_ram_n_23 : std_logic;
  signal gl_ram_n_24, gl_ram_n_25, gl_ram_n_26, gl_ram_n_27, gl_ram_n_28 : std_logic;
  signal gl_ram_n_29, gl_ram_n_30, gl_ram_n_31, gl_ram_n_32, gl_ram_n_33 : std_logic;
  signal gl_ram_n_34, gl_ram_n_35, gl_ram_n_36, gl_ram_n_38, gl_ram_n_40 : std_logic;
  signal gl_ram_n_42, gl_ram_n_44, gl_ram_n_46, gl_ram_n_48, gl_ram_n_50 : std_logic;
  signal gl_ram_n_52, gl_ram_n_54, gl_ram_n_56, gl_ram_n_58, gl_ram_n_60 : std_logic;
  signal gl_ram_n_62, gl_ram_n_64, gl_ram_n_66, gl_ram_n_68, gl_ram_n_70 : std_logic;
  signal gl_ram_n_72, gl_ram_n_74, gl_ram_n_76, gl_ram_n_78, gl_ram_n_80 : std_logic;
  signal gl_ram_n_82, gl_ram_n_84, gl_ram_n_85, gl_ram_n_86, gl_ram_n_87 : std_logic;
  signal gl_ram_n_88, gl_ram_n_89, gl_ram_n_90, gl_ram_n_91, gl_ram_n_92 : std_logic;
  signal gl_ram_n_93, gl_ram_n_94, gl_ram_n_95, gl_ram_n_96, gl_ram_n_97 : std_logic;
  signal gl_ram_n_98, gl_ram_n_99, gl_ram_n_101, gl_ram_n_103, gl_ram_n_105 : std_logic;
  signal gl_ram_n_106, gl_ram_n_107, gl_ram_n_108, gl_ram_n_109, gl_ram_n_110 : std_logic;
  signal gl_ram_n_111, gl_ram_n_112, gl_ram_n_113, gl_ram_n_116, gl_ram_n_118 : std_logic;
  signal gl_ram_n_120, gl_ram_n_121, gl_ram_n_122, gl_ram_n_124, gl_ram_n_125 : std_logic;
  signal gl_ram_n_126, gl_ram_n_127, gl_ram_n_128, gl_ram_n_131, gl_ram_n_132 : std_logic;
  signal gl_ram_n_135, gl_ram_n_137, gl_ram_n_143, gl_ram_n_145, gl_ram_n_146 : std_logic;
  signal gl_ram_n_148, gl_ram_n_150, gl_ram_n_153, gl_ram_n_156, gl_ram_n_157 : std_logic;
  signal gl_ram_n_159, gl_ram_n_161, gl_ram_n_162, gl_ram_n_163, gl_ram_n_164 : std_logic;
  signal gl_ram_n_166, gl_ram_n_168, gl_ram_n_169, gl_ram_n_171, gl_ram_n_173 : std_logic;
  signal gl_ram_n_174, gl_ram_n_176, gl_ram_n_178, gl_ram_n_179, gl_ram_n_181 : std_logic;
  signal gl_ram_n_183, gl_ram_n_185, gl_ram_n_186, gl_ram_n_187, gl_ram_n_188 : std_logic;
  signal gl_ram_n_189, gl_ram_n_191, gl_ram_n_192, gl_ram_n_194, gl_ram_n_201 : std_logic;
  signal gl_ram_n_202, gl_ram_n_203, gl_ram_n_204, gl_ram_n_205, gl_ram_n_207 : std_logic;
  signal gl_ram_n_209, gl_ram_n_213, gl_ram_n_214, gl_ram_n_215, gl_ram_n_216 : std_logic;
  signal gl_ram_n_218, gl_ram_n_220, gl_ram_n_221, gl_ram_n_222, gl_ram_n_224 : std_logic;
  signal gl_ram_n_225, gl_ram_n_226, gl_ram_n_227, gl_ram_n_228, gl_ram_n_229 : std_logic;
  signal gl_ram_n_231, gl_ram_n_232, gl_ram_n_235, gl_ram_n_239, gl_ram_n_240 : std_logic;
  signal gl_ram_n_241, gl_ram_n_242, gl_ram_n_243, gl_ram_n_245, gl_ram_n_246 : std_logic;
  signal gl_ram_n_249, gl_ram_n_251, gl_ram_n_252, gl_ram_n_253, gl_ram_n_254 : std_logic;
  signal gl_ram_n_255, gl_ram_n_256, gl_ram_n_258, gl_ram_n_259, gl_ram_n_260 : std_logic;
  signal gl_ram_n_261, gl_ram_n_263, gl_ram_n_264, gl_ram_n_265, gl_ram_n_267 : std_logic;
  signal gl_ram_n_269, gl_ram_n_270, gl_ram_n_271, gl_ram_n_272, gl_ram_n_273 : std_logic;
  signal gl_ram_n_274, gl_ram_n_276, gl_ram_n_277, gl_ram_n_279, gl_ram_n_281 : std_logic;
  signal gl_ram_n_282, gl_ram_n_283, gl_ram_n_285, gl_ram_n_286, gl_ram_n_288 : std_logic;
  signal gl_ram_n_289, gl_ram_n_290, gl_ram_n_291, gl_ram_n_292, gl_ram_n_293 : std_logic;
  signal gl_ram_n_294, gl_ram_n_296, gl_ram_n_297, gl_ram_n_299, gl_ram_n_300 : std_logic;
  signal gl_ram_n_301, gl_ram_n_303, gl_ram_n_304, gl_ram_n_305, gl_ram_n_307 : std_logic;
  signal gl_ram_n_309, gl_ram_n_310, gl_ram_n_311, gl_ram_n_312, gl_ram_n_315 : std_logic;
  signal gl_ram_n_316, gl_ram_n_322, gl_ram_n_324, gl_ram_n_326, gl_ram_n_330 : std_logic;
  signal gl_ram_n_331, gl_ram_n_332, gl_ram_n_333, gl_ram_n_335, gl_ram_n_336 : std_logic;
  signal gl_ram_n_339, gl_ram_n_340, gl_ram_n_343, gl_ram_n_345, gl_ram_n_346 : std_logic;
  signal gl_ram_n_348, gl_ram_n_350, gl_ram_n_351, gl_ram_n_353, gl_ram_n_354 : std_logic;
  signal gl_ram_n_357, gl_ram_n_359, gl_ram_n_360, gl_ram_n_361, gl_ram_n_362 : std_logic;
  signal gl_ram_n_366, gl_ram_n_371, gl_ram_n_373, gl_ram_n_378, gl_ram_n_379 : std_logic;
  signal gl_ram_n_380, gl_ram_n_381, gl_ram_n_387, gl_ram_n_388, gl_ram_n_389 : std_logic;
  signal gl_ram_n_390, gl_ram_n_391, gl_ram_n_393, gl_ram_n_394, gl_ram_n_395 : std_logic;
  signal gl_ram_n_396, gl_ram_n_398, gl_ram_n_399, gl_ram_n_400, gl_ram_n_401 : std_logic;
  signal gl_ram_n_403, gl_ram_n_404, gl_ram_n_405, gl_ram_n_406, gl_ram_n_407 : std_logic;
  signal gl_ram_n_408, gl_ram_n_409, gl_ram_n_410, gl_ram_n_414, gl_ram_n_415 : std_logic;
  signal gl_ram_n_417, gl_ram_n_424, gl_ram_n_426, gl_ram_n_433, gl_ram_n_439 : std_logic;
  signal gl_ram_n_450, gl_ram_n_451, gl_ram_n_457, gl_ram_n_458, gl_ram_n_459 : std_logic;
  signal gl_ram_n_463, gl_ram_n_465, gl_ram_n_467, gl_ram_n_471, gl_ram_n_472 : std_logic;
  signal gl_ram_n_475, gl_ram_n_481, gl_ram_n_482, gl_ram_n_484, gl_ram_n_485 : std_logic;
  signal gl_ram_n_492, gl_ram_n_495, gl_ram_n_496, gl_ram_n_498, gl_ram_n_499 : std_logic;
  signal gl_ram_n_500, gl_ram_n_503, gl_ram_n_507, gl_ram_n_508, gl_ram_n_510 : std_logic;
  signal gl_ram_n_517, gl_ram_n_518, gl_ram_n_526, gl_ram_n_541, gl_ram_n_543 : std_logic;
  signal gl_ram_n_545, gl_ram_n_547, gl_ram_n_548, gl_ram_n_550, gl_ram_n_552 : std_logic;
  signal gl_ram_n_553, gl_ram_n_554, gl_ram_n_555, gl_ram_n_556, gl_ram_n_557 : std_logic;
  signal gl_ram_n_558, gl_ram_n_559, gl_ram_n_560, gl_ram_n_561, gl_ram_n_562 : std_logic;
  signal gl_ram_n_563, gl_ram_n_564, gl_ram_n_565, gl_ram_n_567, gl_ram_n_568 : std_logic;
  signal gl_ram_n_570, gl_ram_n_571, gl_ram_n_572, gl_ram_n_573, gl_ram_n_575 : std_logic;
  signal gl_ram_n_576, gl_ram_n_577, gl_ram_n_578, gl_ram_n_579, gl_ram_n_580 : std_logic;
  signal gl_ram_n_581, gl_ram_n_582, gl_ram_n_583, gl_ram_n_584, gl_ram_n_585 : std_logic;
  signal gl_ram_n_586, gl_ram_n_587, gl_ram_n_588, gl_ram_n_589, gl_ram_n_590 : std_logic;
  signal gl_ram_n_591, gl_ram_n_592, gl_ram_n_593, gl_ram_n_594, gl_ram_n_595 : std_logic;
  signal gl_ram_n_596, gl_ram_n_597, gl_ram_n_599, gl_ram_n_600, gl_ram_n_601 : std_logic;
  signal gl_ram_n_602, gl_ram_n_603, gl_ram_n_604, gl_ram_n_605, gl_ram_n_606 : std_logic;
  signal gl_ram_n_607, gl_ram_n_608, gl_ram_n_609, gl_ram_n_610, gl_ram_n_611 : std_logic;
  signal gl_ram_n_613, gl_ram_n_614, gl_ram_n_615, gl_ram_n_616, gl_ram_n_617 : std_logic;
  signal gl_ram_n_618, gl_ram_n_619, gl_ram_n_620, gl_ram_n_621, gl_ram_n_622 : std_logic;
  signal gl_ram_n_623, gl_ram_n_624, gl_ram_n_625, gl_ram_n_626, gl_ram_n_627 : std_logic;
  signal gl_ram_n_628, gl_ram_n_629, gl_ram_n_630, gl_ram_n_631, gl_ram_n_632 : std_logic;
  signal gl_ram_n_633, gl_ram_n_634, gl_ram_n_635, gl_ram_n_636, gl_ram_n_637 : std_logic;
  signal gl_ram_n_638, gl_ram_n_639, gl_ram_n_640, gl_ram_n_641, gl_ram_n_642 : std_logic;
  signal gl_ram_n_643, gl_ram_n_644, gl_ram_n_645, gl_ram_n_646, gl_ram_n_647 : std_logic;
  signal gl_ram_n_648, gl_ram_n_649, gl_ram_n_650, gl_ram_n_651, gl_ram_n_652 : std_logic;
  signal gl_ram_n_653, gl_ram_n_657, gl_ram_n_658, gl_ram_n_659, gl_ram_n_660 : std_logic;
  signal gl_ram_n_661, gl_ram_n_662, gl_ram_n_663, gl_ram_n_664, gl_ram_n_665 : std_logic;
  signal gl_ram_n_668, gl_ram_n_669, gl_ram_n_671, gl_ram_n_672, gl_ram_n_673 : std_logic;
  signal gl_ram_n_674, gl_ram_n_675, gl_ram_n_676, gl_ram_n_677, gl_ram_n_678 : std_logic;
  signal gl_ram_n_679, gl_ram_n_680, gl_ram_n_681, gl_ram_n_682, gl_ram_n_683 : std_logic;
  signal gl_ram_n_684, gl_ram_n_685, gl_ram_n_686, gl_ram_n_687, gl_ram_n_688 : std_logic;
  signal gl_ram_n_689, gl_ram_n_690, gl_ram_n_691, gl_ram_n_692, gl_ram_n_693 : std_logic;
  signal gl_ram_n_694, gl_ram_n_695, gl_ram_n_696, gl_ram_n_697, gl_ram_n_698 : std_logic;
  signal gl_ram_n_699, gl_ram_n_700, gl_ram_n_701, gl_ram_n_702, gl_ram_n_703 : std_logic;
  signal gl_ram_n_704, gl_ram_n_705, gl_ram_n_706, gl_ram_n_707, gl_ram_n_708 : std_logic;
  signal gl_ram_n_709, gl_ram_n_710, gl_ram_n_711, gl_ram_n_712, gl_ram_n_713 : std_logic;
  signal gl_ram_n_714, gl_ram_n_715, gl_ram_n_716, gl_ram_n_717, gl_ram_n_718 : std_logic;
  signal gl_ram_n_719, gl_ram_n_720, gl_ram_n_721, gl_ram_n_722, gl_ram_n_723 : std_logic;
  signal gl_ram_n_724, gl_ram_n_725, gl_ram_n_726, gl_ram_n_727, gl_ram_n_728 : std_logic;
  signal gl_ram_n_729, gl_ram_n_730, gl_ram_n_731, gl_ram_n_732, gl_ram_n_733 : std_logic;
  signal gl_ram_n_735, gl_ram_n_736, gl_ram_n_739, gl_ram_n_740, gl_ram_n_741 : std_logic;
  signal gl_ram_n_742, gl_ram_n_743, gl_ram_n_744, gl_ram_n_745, gl_ram_n_746 : std_logic;
  signal gl_ram_n_747, gl_ram_n_748, gl_ram_n_749, gl_ram_n_750, gl_ram_n_751 : std_logic;
  signal gl_ram_n_752, gl_ram_n_753, gl_ram_n_754, gl_ram_n_755, gl_ram_n_756 : std_logic;
  signal gl_ram_n_757, gl_ram_n_758, gl_ram_n_759, gl_ram_n_760, gl_ram_n_761 : std_logic;
  signal gl_ram_n_762, gl_ram_n_763, gl_ram_n_764, gl_ram_n_765, gl_ram_n_766 : std_logic;
  signal gl_ram_n_767, gl_ram_n_768, gl_ram_n_769, gl_ram_n_770, gl_ram_n_771 : std_logic;
  signal gl_ram_n_772, gl_ram_n_773, gl_ram_n_774, gl_ram_n_775, gl_ram_n_776 : std_logic;
  signal gl_ram_n_777, gl_ram_n_778, gl_ram_n_779, gl_ram_n_780, gl_ram_n_781 : std_logic;
  signal gl_ram_n_782, gl_ram_n_783, gl_ram_n_784, gl_ram_n_785, gl_ram_n_786 : std_logic;
  signal gl_ram_n_787, gl_ram_n_788, gl_ram_n_789, gl_ram_n_790, gl_ram_n_791 : std_logic;
  signal gl_ram_n_792, gl_ram_n_793, gl_ram_n_794, gl_ram_n_795, gl_ram_n_796 : std_logic;
  signal gl_ram_n_797, gl_ram_n_798, gl_ram_n_799, gl_ram_n_800, gl_ram_n_801 : std_logic;
  signal gl_ram_n_802, gl_ram_n_803, gl_ram_n_804, gl_ram_n_805, gl_ram_n_806 : std_logic;
  signal gl_ram_n_807, gl_ram_n_808, gl_ram_n_809, gl_ram_n_810, gl_ram_n_811 : std_logic;
  signal gl_ram_n_812, gl_ram_n_813, gl_ram_n_814, gl_ram_n_815, gl_ram_n_816 : std_logic;
  signal gl_ram_n_817, gl_ram_n_818, gl_ram_n_819, gl_ram_n_820, gl_ram_n_821 : std_logic;
  signal gl_ram_n_822, gl_ram_n_823, gl_ram_n_824, gl_ram_n_825, gl_ram_n_826 : std_logic;
  signal gl_ram_n_827, gl_ram_n_828, gl_ram_n_829, gl_ram_n_830, gl_ram_n_831 : std_logic;
  signal gl_ram_n_832, gl_ram_n_833, gl_ram_n_834, gl_ram_n_835, gl_ram_n_836 : std_logic;
  signal gl_ram_n_837, gl_ram_n_838, gl_ram_n_839, gl_ram_n_840, gl_ram_n_841 : std_logic;
  signal gl_ram_n_842, gl_ram_n_843, gl_ram_n_844, gl_ram_n_845, gl_ram_n_846 : std_logic;
  signal gl_ram_n_847, gl_ram_n_848, gl_ram_n_849, gl_ram_n_850, gl_ram_n_851 : std_logic;
  signal gl_ram_n_852, gl_ram_n_853, gl_ram_n_854, gl_ram_n_855, gl_ram_n_856 : std_logic;
  signal gl_ram_n_857, gl_ram_n_858, gl_ram_n_859, gl_ram_n_860, gl_ram_n_861 : std_logic;
  signal gl_ram_n_862, gl_ram_n_863, gl_ram_n_864, gl_ram_n_865, gl_ram_n_866 : std_logic;
  signal gl_ram_n_867, gl_ram_n_868, gl_ram_n_869, gl_ram_n_870, gl_ram_n_871 : std_logic;
  signal gl_ram_n_872, gl_ram_n_873, gl_ram_n_874, gl_ram_n_875, gl_ram_n_876 : std_logic;
  signal gl_ram_n_877, gl_ram_n_878, gl_ram_n_879, gl_ram_n_880, gl_ram_n_881 : std_logic;
  signal gl_ram_n_882, gl_ram_n_883, gl_ram_n_884, gl_ram_n_885, gl_ram_n_886 : std_logic;
  signal gl_ram_n_887, gl_ram_n_888, gl_ram_n_889, gl_ram_n_890, gl_ram_n_891 : std_logic;
  signal gl_ram_n_892, gl_ram_n_893, gl_ram_n_894, gl_ram_n_895, gl_ram_n_896 : std_logic;
  signal gl_ram_n_897, gl_ram_n_898, gl_ram_n_899, gl_ram_n_900, gl_ram_n_901 : std_logic;
  signal gl_ram_n_902, gl_ram_n_903, gl_ram_n_904, gl_ram_n_905, gl_ram_n_906 : std_logic;
  signal gl_ram_n_907, gl_ram_n_908, gl_ram_n_909, gl_ram_n_910, gl_ram_n_911 : std_logic;
  signal gl_ram_n_912, gl_ram_n_913, gl_ram_n_914, gl_ram_n_915, gl_ram_n_916 : std_logic;
  signal gl_ram_n_917, gl_ram_n_918, gl_ram_n_919, gl_ram_n_920, gl_ram_n_921 : std_logic;
  signal gl_ram_n_922, gl_ram_n_923, gl_ram_n_924, gl_ram_n_925, gl_ram_n_926 : std_logic;
  signal gl_ram_n_927, gl_ram_n_928, gl_ram_n_929, gl_ram_n_930, gl_ram_n_931 : std_logic;
  signal gl_ram_n_932, gl_ram_n_933, gl_ram_n_934, gl_ram_n_935, gl_ram_n_936 : std_logic;
  signal gl_ram_n_937, gl_ram_n_938, gl_ram_n_939, gl_ram_n_940, gl_ram_n_941 : std_logic;
  signal gl_ram_n_942, gl_ram_n_943, gl_ram_n_944, gl_ram_n_945, gl_ram_n_946 : std_logic;
  signal gl_ram_n_947, gl_ram_n_948, gl_ram_n_949, gl_ram_n_950, gl_ram_n_951 : std_logic;
  signal gl_ram_n_952, gl_ram_n_953, gl_ram_n_954, gl_ram_n_955, gl_ram_n_956 : std_logic;
  signal gl_ram_n_957, gl_ram_n_958, gl_ram_n_959, gl_ram_n_960, gl_ram_n_961 : std_logic;
  signal gl_ram_n_962, gl_ram_n_963, gl_ram_n_964, gl_ram_n_965, gl_ram_n_966 : std_logic;
  signal gl_ram_n_967, gl_ram_n_968, gl_ram_n_969, gl_ram_n_970, gl_ram_n_971 : std_logic;
  signal gl_ram_n_972, gl_ram_n_973, gl_ram_n_974, gl_ram_n_975, gl_ram_n_976 : std_logic;
  signal gl_ram_n_977, gl_ram_n_978, gl_ram_n_979, gl_ram_n_980, gl_ram_n_981 : std_logic;
  signal gl_ram_n_982, gl_ram_n_983, gl_ram_n_984, gl_ram_n_985, gl_ram_n_986 : std_logic;
  signal gl_ram_n_987, gl_ram_n_988, gl_ram_n_989, gl_ram_n_990, gl_ram_n_991 : std_logic;
  signal gl_ram_n_992, gl_ram_n_993, gl_ram_n_994, gl_ram_n_995, gl_ram_n_996 : std_logic;
  signal gl_ram_n_997, gl_ram_n_998, gl_ram_n_999, gl_ram_n_1000, gl_ram_n_1001 : std_logic;
  signal gl_ram_n_1002, gl_ram_n_1003, gl_ram_n_1004, gl_ram_n_1005, gl_ram_n_1006 : std_logic;
  signal gl_ram_n_1007, gl_ram_n_1008, gl_ram_n_1009, gl_ram_n_1010, gl_ram_n_1011 : std_logic;
  signal gl_ram_n_1012, gl_ram_n_1013, gl_ram_n_1014, gl_ram_n_1015, gl_ram_n_1016 : std_logic;
  signal gl_ram_n_1017, gl_ram_n_1018, gl_ram_n_1019, gl_ram_n_1020, gl_ram_n_1021 : std_logic;
  signal gl_ram_n_1022, gl_ram_n_1023, gl_ram_n_1024, gl_ram_n_1025, gl_ram_n_1026 : std_logic;
  signal gl_ram_n_1027, gl_ram_n_1028, gl_ram_n_1029, gl_ram_n_1030, gl_ram_n_1031 : std_logic;
  signal gl_ram_n_1032, gl_ram_n_1033, gl_ram_n_1034, gl_ram_n_1035, gl_ram_n_1036 : std_logic;
  signal gl_ram_n_1037, gl_ram_n_1038, gl_ram_n_1039, gl_ram_n_1040, gl_ram_n_1041 : std_logic;
  signal gl_ram_n_1042, gl_ram_n_1043, gl_ram_n_1044, gl_ram_n_1045, gl_ram_n_1046 : std_logic;
  signal gl_ram_n_1047, gl_ram_n_1048, gl_ram_n_1049, gl_ram_n_1050, gl_ram_n_1051 : std_logic;
  signal gl_ram_n_1052, gl_ram_n_1053, gl_ram_n_1054, gl_ram_n_1055, gl_ram_n_1056 : std_logic;
  signal gl_ram_n_1057, gl_ram_n_1058, gl_ram_n_1059, gl_ram_n_1060, gl_ram_n_1061 : std_logic;
  signal gl_ram_n_1062, gl_ram_n_1063, gl_ram_n_1064, gl_ram_n_1065, gl_ram_n_1066 : std_logic;
  signal gl_ram_n_1067, gl_ram_n_1068, gl_ram_n_1069, gl_ram_n_1070, gl_ram_n_1071 : std_logic;
  signal gl_ram_n_1072, gl_ram_n_1073, gl_ram_n_1074, gl_ram_n_1075, gl_ram_n_1076 : std_logic;
  signal gl_ram_n_1077, gl_ram_n_1078, gl_ram_n_1079, gl_ram_n_1080, gl_ram_n_1081 : std_logic;
  signal gl_ram_n_1082, gl_ram_n_1083, gl_ram_n_1084, gl_ram_n_1085, gl_ram_n_1086 : std_logic;
  signal gl_ram_n_1087, gl_ram_n_1088, gl_ram_n_1089, gl_ram_n_1090, gl_ram_n_1091 : std_logic;
  signal gl_ram_n_1092, gl_ram_n_1093, gl_ram_n_1094, gl_ram_n_1095, gl_ram_n_1096 : std_logic;
  signal gl_ram_n_1097, gl_ram_n_1098, gl_ram_n_1099, gl_ram_n_1100, gl_ram_n_1101 : std_logic;
  signal gl_ram_n_1102, gl_ram_n_1103, gl_ram_n_1104, gl_ram_n_1105, gl_ram_n_1106 : std_logic;
  signal gl_ram_n_1107, gl_ram_n_1108, gl_ram_n_1109, gl_ram_n_1110, gl_ram_n_1111 : std_logic;
  signal gl_ram_n_1112, gl_ram_n_1114, gl_ram_n_1116, gl_ram_n_1118, gl_ram_n_1120 : std_logic;
  signal gl_ram_n_1122, gl_ram_n_1124, gl_ram_n_1126, gl_ram_n_1128, gl_ram_n_1130 : std_logic;
  signal gl_ram_n_1132, gl_ram_n_1134, gl_ram_n_1136, gl_ram_n_1138, gl_ram_n_1140 : std_logic;
  signal gl_ram_n_1142, gl_ram_n_1144, gl_ram_n_1146, gl_ram_n_1148, gl_ram_n_1150 : std_logic;
  signal gl_ram_n_1152, gl_ram_n_1154, gl_ram_n_1156, gl_ram_n_1158, gl_ram_n_1160 : std_logic;
  signal gl_ram_n_1162, gl_ram_n_1164, gl_ram_n_1166, gl_ram_n_1168, gl_ram_n_1170 : std_logic;
  signal gl_ram_n_1172, gl_ram_n_1174, gl_ram_n_1176, gl_ram_n_1178, gl_ram_n_1180 : std_logic;
  signal gl_ram_n_1182, gl_ram_n_1184, gl_ram_n_1186, gl_ram_n_1188, gl_ram_n_1190 : std_logic;
  signal gl_ram_n_1192, gl_ram_n_1194, gl_ram_n_1196, gl_ram_n_1198, gl_ram_n_1200 : std_logic;
  signal gl_ram_n_1202, gl_ram_n_1204, gl_ram_n_1206, gl_ram_n_1208, gl_ram_n_1210 : std_logic;
  signal gl_ram_n_1212, gl_ram_n_1214, gl_ram_n_1216, gl_ram_n_1218, gl_ram_n_1220 : std_logic;
  signal gl_ram_n_1222, gl_ram_n_1224, gl_ram_n_1226, gl_ram_n_1228, gl_ram_n_1230 : std_logic;
  signal gl_ram_n_1232, gl_ram_n_1234, gl_ram_n_1236, gl_ram_n_1238, gl_ram_n_1240 : std_logic;
  signal gl_ram_n_1242, gl_ram_n_1244, gl_ram_n_1246, gl_ram_n_1248, gl_ram_n_1250 : std_logic;
  signal gl_ram_n_1252, gl_ram_n_1254, gl_ram_n_1256, gl_ram_n_1258, gl_ram_n_1260 : std_logic;
  signal gl_ram_n_1262, gl_ram_n_1264, gl_ram_n_1266, gl_ram_n_1268, gl_ram_n_1270 : std_logic;
  signal gl_ram_n_1272, gl_ram_n_1274, gl_ram_n_1276, gl_ram_n_1278, gl_ram_n_1280 : std_logic;
  signal gl_ram_n_1282, gl_ram_n_1284, gl_ram_n_1286, gl_ram_n_1288, gl_ram_n_1290 : std_logic;
  signal gl_ram_n_1292, gl_ram_n_1294, gl_ram_n_1296, gl_ram_n_1298, gl_ram_n_1300 : std_logic;
  signal gl_ram_n_1302, gl_ram_n_1304, gl_ram_n_1306, gl_ram_n_1308, gl_ram_n_1310 : std_logic;
  signal gl_ram_n_1311, gl_ram_n_1320, gl_ram_n_1436, gl_ram_n_1437, gl_ram_n_1438 : std_logic;
  signal gl_ram_n_1439, gl_ram_n_1440, gl_ram_n_1444, gl_ram_n_1445, gl_ram_n_1446 : std_logic;
  signal gl_ram_n_1447, gl_ram_n_1448, gl_ram_n_1449, gl_ram_n_1450, gl_ram_n_1451 : std_logic;
  signal gl_ram_n_1452, gl_ram_n_1453, gl_ram_n_1454, gl_ram_n_1455, gl_ram_n_1456 : std_logic;
  signal gl_ram_n_1457, gl_ram_n_1458, gl_ram_n_1459, gl_ram_n_1460, gl_ram_n_1461 : std_logic;
  signal gl_ram_n_1462, gl_ram_n_1463, gl_ram_n_1464, gl_ram_n_1465, gl_ram_n_1466 : std_logic;
  signal gl_ram_n_1467, gl_ram_n_1468, gl_ram_n_1469, gl_ram_n_1470, gl_ram_n_1471 : std_logic;
  signal gl_ram_n_1472, gl_ram_n_1473, gl_ram_n_1474, gl_ram_n_1475, gl_ram_n_1476 : std_logic;
  signal gl_ram_n_1477, gl_ram_n_1478, gl_ram_n_1479, gl_ram_n_1480, gl_ram_n_1481 : std_logic;
  signal gl_ram_n_1482, gl_ram_n_1483, gl_ram_n_1484, gl_ram_n_1485, gl_ram_n_1486 : std_logic;
  signal gl_ram_n_1487, gl_ram_n_1488, gl_ram_n_1489, gl_ram_n_1490, gl_ram_n_1491 : std_logic;
  signal gl_ram_n_1492, gl_ram_n_1493, gl_ram_n_1494, gl_ram_n_1495, gl_ram_n_1496 : std_logic;
  signal gl_ram_n_1497, gl_ram_n_1498, gl_ram_n_1499, gl_ram_n_1500, gl_ram_n_1501 : std_logic;
  signal gl_ram_n_1502, gl_ram_n_1503, gl_ram_n_1504, gl_ram_n_1505, gl_ram_n_1506 : std_logic;
  signal gl_ram_n_1507, gl_ram_n_1508, gl_ram_n_1509, gl_ram_n_1510, gl_ram_n_1511 : std_logic;
  signal gl_ram_n_1512, gl_ram_n_1513, gl_ram_n_1514, gl_ram_n_1515, gl_ram_n_1516 : std_logic;
  signal gl_ram_n_1517, gl_ram_n_1518, gl_ram_n_1519, gl_ram_n_1520, gl_ram_n_1521 : std_logic;
  signal gl_ram_n_1522, gl_ram_n_1523, gl_ram_n_1524, gl_ram_n_1525, gl_ram_n_1526 : std_logic;
  signal gl_ram_n_1527, gl_ram_n_1528, gl_ram_n_1529, gl_ram_n_1530, gl_ram_n_1531 : std_logic;
  signal gl_ram_n_1532, gl_ram_n_1533, gl_ram_n_1534, gl_ram_n_1535, gl_ram_n_1536 : std_logic;
  signal gl_ram_n_1537, gl_ram_n_1538, gl_ram_n_1539, gl_ram_n_1540, gl_ram_n_1541 : std_logic;
  signal gl_ram_n_1542, gl_ram_n_1543, gl_ram_n_1544, gl_ram_n_1545, gl_ram_n_1546 : std_logic;
  signal gl_ram_n_1547, gl_ram_n_1548, gl_ram_n_1549, gl_ram_n_1550, gl_ram_n_1551 : std_logic;
  signal gl_ram_n_1552, gl_rom_n_0, gl_rom_n_1, gl_rom_n_2, gl_rom_n_3 : std_logic;
  signal gl_rom_n_4, gl_rom_n_5, gl_rom_n_6, gl_rom_n_7, gl_rom_n_8 : std_logic;
  signal gl_rom_n_9, gl_rom_n_10, gl_rom_n_11, gl_rom_n_12, gl_rom_n_13 : std_logic;
  signal gl_rom_n_14, gl_rom_n_15, gl_rom_n_16, gl_rom_n_17, gl_rom_n_18 : std_logic;
  signal gl_rom_n_19, gl_rom_n_20, gl_rom_n_21, gl_rom_n_22, gl_rom_n_23 : std_logic;
  signal gl_rom_n_24, gl_rom_n_25, gl_rom_n_26, gl_rom_n_27, gl_rom_n_28 : std_logic;
  signal gl_rom_n_29, gl_rom_n_30, gl_rom_n_31, gl_rom_n_32, gl_rom_n_33 : std_logic;
  signal gl_rom_n_34, gl_rom_n_35, gl_rom_n_36, gl_rom_n_37, gl_rom_n_38 : std_logic;
  signal gl_rom_n_39, gl_rom_n_40, gl_rom_n_41, gl_rom_n_42, gl_rom_n_43 : std_logic;
  signal gl_rom_n_44, gl_rom_n_45, gl_rom_n_46, gl_rom_n_47, gl_rom_n_48 : std_logic;
  signal gl_rom_n_49, gl_rom_n_50, gl_rom_n_51, gl_rom_n_52, gl_rom_n_53 : std_logic;
  signal gl_rom_n_54, gl_rom_n_55, gl_rom_n_56, gl_rom_n_57, gl_rom_n_58 : std_logic;
  signal gl_rom_n_59, gl_rom_n_60, gl_rom_n_61, gl_rom_n_62, gl_rom_n_63 : std_logic;
  signal gl_rom_n_64, gl_rom_n_65, gl_rom_n_66, gl_rom_n_67, gl_rom_n_68 : std_logic;
  signal gl_rom_n_69, gl_rom_n_70, gl_rom_n_71, gl_rom_n_72, gl_rom_n_73 : std_logic;
  signal gl_rom_n_74, gl_rom_n_75, gl_rom_n_76, gl_rom_n_77, gl_rom_n_78 : std_logic;
  signal gl_rom_n_79, gl_rom_n_80, gl_rom_n_81, gl_rom_n_82, gl_rom_n_83 : std_logic;
  signal gl_rom_n_84, gl_rom_n_85, gl_rom_n_86, gl_rom_n_87, gl_rom_n_88 : std_logic;
  signal gl_rom_n_89, gl_rom_n_90, gl_rom_n_91, gl_rom_n_92, gl_rom_n_93 : std_logic;
  signal gl_rom_n_94, gl_rom_n_95, gl_rom_n_96, gl_rom_n_97, gl_rom_n_98 : std_logic;
  signal gl_rom_n_99, gl_rom_n_100, gl_rom_n_101, gl_rom_n_102, gl_rom_n_103 : std_logic;
  signal gl_rom_n_104, gl_rom_n_105, gl_rom_n_106, gl_rom_n_107, gl_rom_n_108 : std_logic;
  signal gl_rom_n_109, gl_rom_n_110, gl_rom_n_111, gl_rom_n_112, gl_rom_n_113 : std_logic;
  signal gl_rom_n_114, gl_rom_n_115, gl_rom_n_116, gl_rom_n_117, gl_rom_n_118 : std_logic;
  signal gl_rom_n_119, gl_rom_n_120, gl_rom_n_121, gl_rom_n_122, gl_rom_n_123 : std_logic;
  signal gl_rom_n_124, gl_rom_n_125, gl_rom_n_126, gl_rom_n_127, gl_rom_n_128 : std_logic;
  signal gl_rom_n_129, gl_rom_n_130, gl_rom_n_131, gl_rom_n_132, gl_rom_n_133 : std_logic;
  signal gl_rom_n_134, gl_rom_n_135, gl_rom_n_136, gl_rom_n_137, gl_rom_n_138 : std_logic;
  signal gl_rom_n_139, gl_rom_n_140, gl_rom_n_141, gl_rom_n_142, gl_rom_n_143 : std_logic;
  signal gl_rom_n_144, gl_rom_n_145, gl_rom_n_146, gl_rom_n_147, gl_rom_n_148 : std_logic;
  signal gl_rom_n_149, gl_rom_n_150, gl_rom_n_151, gl_rom_n_152, gl_rom_n_153 : std_logic;
  signal gl_rom_n_154, gl_rom_n_155, gl_rom_n_156, gl_rom_n_157, gl_rom_n_158 : std_logic;
  signal gl_rom_n_159, gl_rom_n_160, gl_rom_n_161, gl_rom_n_162, gl_rom_n_163 : std_logic;
  signal gl_rom_n_164, gl_rom_n_165, gl_rom_n_166, gl_rom_n_167, gl_rom_n_168 : std_logic;
  signal gl_rom_n_169, gl_rom_n_170, gl_rom_n_171, gl_rom_n_172, gl_rom_n_173 : std_logic;
  signal gl_rom_n_174, gl_rom_n_175, gl_rom_n_176, gl_rom_n_177, gl_rom_n_178 : std_logic;
  signal gl_rom_n_179, gl_rom_n_180, gl_rom_n_181, gl_rom_n_182, gl_rom_n_183 : std_logic;
  signal gl_rom_n_184, gl_rom_n_185, gl_rom_n_186, gl_rom_n_187, gl_rom_n_188 : std_logic;
  signal gl_rom_n_189, gl_rom_n_190, gl_rom_n_191, gl_rom_n_192, gl_rom_n_193 : std_logic;
  signal gl_rom_n_194, gl_rom_n_195, gl_rom_n_196, gl_rom_n_197, gl_rom_n_198 : std_logic;
  signal gl_rom_n_199, gl_rom_n_200, gl_rom_n_201, gl_rom_n_202, gl_rom_n_203 : std_logic;
  signal gl_rom_n_204, gl_rom_n_205, gl_rom_n_206, gl_rom_n_207, gl_rom_n_208 : std_logic;
  signal gl_rom_n_209, gl_rom_n_210, gl_rom_n_211, gl_rom_n_212, gl_rom_n_213 : std_logic;
  signal gl_rom_n_214, gl_rom_n_215, gl_rom_n_216, gl_rom_n_217, gl_rom_n_218 : std_logic;
  signal gl_rom_n_219, gl_rom_n_220, gl_rom_n_221, gl_rom_n_222, gl_rom_n_223 : std_logic;
  signal gl_rom_n_224, gl_rom_n_225, gl_rom_n_226, gl_rom_n_227, gl_rom_n_228 : std_logic;
  signal gl_rom_n_229, gl_rom_n_230, gl_rom_n_231, gl_rom_n_232, gl_rom_n_233 : std_logic;
  signal gl_rom_n_234, gl_rom_n_235, gl_rom_n_236, gl_rom_n_237, gl_rom_n_238 : std_logic;
  signal gl_rom_n_239, gl_rom_n_240, gl_rom_n_241, gl_rom_n_242, gl_rom_n_243 : std_logic;
  signal gl_rom_n_244, gl_rom_n_245, gl_rom_n_246, gl_rom_n_247, gl_rom_n_248 : std_logic;
  signal gl_rom_n_249, gl_rom_n_250, gl_rom_n_251, gl_rom_n_252, gl_rom_n_253 : std_logic;
  signal gl_rom_n_254, gl_rom_n_255, gl_rom_n_256, gl_rom_n_257, gl_rom_n_258 : std_logic;
  signal gl_rom_n_259, gl_rom_n_260, gl_rom_n_261, gl_rom_n_262, gl_rom_n_263 : std_logic;
  signal gl_rom_n_264, gl_rom_n_265, gl_rom_n_266, gl_rom_n_267, gl_rom_n_268 : std_logic;
  signal gl_rom_n_269, gl_rom_n_270, gl_rom_n_271, gl_rom_n_272, gl_rom_n_273 : std_logic;
  signal gl_rom_n_274, gl_rom_n_275, gl_rom_n_276, gl_rom_n_277, gl_rom_n_278 : std_logic;
  signal gl_rom_n_279, gl_rom_n_280, gl_rom_n_281, gl_rom_n_282, gl_rom_n_283 : std_logic;
  signal gl_rom_n_284, gl_rom_n_285, gl_rom_n_286, gl_rom_n_287, gl_rom_n_288 : std_logic;
  signal gl_rom_n_289, gl_rom_n_290, gl_rom_n_291, gl_rom_n_292, gl_rom_n_293 : std_logic;
  signal gl_rom_n_294, gl_rom_n_295, gl_rom_n_296, gl_rom_n_297, gl_rom_n_298 : std_logic;
  signal gl_rom_n_299, gl_rom_n_300, gl_rom_n_301, gl_rom_n_302, gl_rom_n_303 : std_logic;
  signal gl_rom_n_304, gl_rom_n_305, gl_rom_n_306, gl_rom_n_307, gl_rom_n_308 : std_logic;
  signal gl_rom_n_309, gl_rom_n_310, gl_rom_n_311, gl_rom_n_312, gl_rom_n_313 : std_logic;
  signal gl_rom_n_314, gl_rom_n_315, gl_rom_n_316, gl_rom_n_317, gl_rom_n_318 : std_logic;
  signal gl_rom_n_319, gl_rom_n_320, gl_rom_n_321, gl_rom_n_322, gl_rom_n_323 : std_logic;
  signal gl_rom_n_324, gl_rom_n_325, gl_rom_n_326, gl_rom_n_327, gl_rom_n_328 : std_logic;
  signal gl_rom_n_329, gl_rom_n_330, gl_rom_n_331, gl_rom_n_332, gl_rom_n_333 : std_logic;
  signal gl_rom_n_334, gl_rom_n_335, gl_rom_n_336, gl_rom_n_337, gl_rom_n_338 : std_logic;
  signal gl_rom_n_339, gl_rom_n_340, gl_rom_n_341, gl_rom_n_342, gl_rom_n_343 : std_logic;
  signal gl_rom_n_344, gl_rom_n_345, gl_rom_n_346, gl_rom_n_347, gl_rom_n_348 : std_logic;
  signal gl_rom_n_349, gl_rom_n_350, gl_rom_n_351, gl_rom_n_352, gl_rom_n_353 : std_logic;
  signal gl_rom_n_354, gl_rom_n_355, gl_rom_n_356, gl_rom_n_357, gl_rom_n_358 : std_logic;
  signal gl_rom_n_359, gl_rom_n_360, gl_rom_n_361, gl_rom_n_362, gl_rom_n_363 : std_logic;
  signal gl_rom_n_364, gl_rom_n_365, gl_rom_n_366, gl_rom_n_367, gl_rom_n_368 : std_logic;
  signal gl_rom_n_369, gl_rom_n_370, gl_rom_n_371, gl_rom_n_372, gl_rom_n_373 : std_logic;
  signal gl_rom_n_374, gl_rom_n_375, gl_rom_n_376, gl_rom_n_377, gl_rom_n_378 : std_logic;
  signal gl_rom_n_379, gl_rom_n_380, gl_rom_n_381, gl_rom_n_382, gl_rom_n_383 : std_logic;
  signal gl_rom_n_384, gl_rom_n_385, gl_rom_n_386, gl_rom_n_387, gl_rom_n_388 : std_logic;
  signal gl_rom_n_389, gl_rom_n_390, gl_rom_n_391, gl_rom_n_392, gl_rom_n_393 : std_logic;
  signal gl_rom_n_394, gl_rom_n_395, gl_rom_n_396, gl_rom_n_397, gl_rom_n_398 : std_logic;
  signal gl_rom_n_399, gl_rom_n_400, gl_rom_n_401, gl_rom_n_402, gl_rom_n_403 : std_logic;
  signal gl_rom_n_404, gl_rom_n_405, gl_rom_n_406, gl_rom_n_407, gl_rom_n_408 : std_logic;
  signal gl_rom_n_409, gl_rom_n_410, gl_rom_n_411, gl_rom_n_412, gl_rom_n_413 : std_logic;
  signal gl_rom_n_414, gl_rom_n_415, gl_rom_n_416, gl_rom_n_417, gl_rom_n_418 : std_logic;
  signal gl_rom_n_419, gl_rom_n_420, gl_rom_n_421, gl_rom_n_422, gl_rom_n_423 : std_logic;
  signal gl_rom_n_424, gl_rom_n_425, gl_rom_n_426, gl_rom_n_427, gl_rom_n_428 : std_logic;
  signal gl_rom_n_429, gl_rom_n_430, gl_rom_n_431, gl_rom_n_432, gl_rom_n_433 : std_logic;
  signal gl_rom_n_434, gl_rom_n_435, gl_rom_n_436, gl_rom_n_437, gl_rom_n_438 : std_logic;
  signal gl_rom_n_439, gl_rom_n_440, gl_rom_n_441, gl_rom_n_442, gl_rom_n_443 : std_logic;
  signal gl_rom_n_444, gl_rom_n_445, gl_rom_n_446, gl_rom_n_447, gl_rom_n_448 : std_logic;
  signal gl_rom_n_449, gl_rom_n_450, gl_rom_n_451, gl_rom_n_452, gl_rom_n_453 : std_logic;
  signal gl_rom_n_454, gl_rom_n_455, gl_rom_n_456, gl_rom_n_457, gl_rom_n_458 : std_logic;
  signal gl_rom_n_459, gl_rom_n_460, gl_rom_n_461, gl_rom_n_462, gl_rom_n_463 : std_logic;
  signal gl_rom_n_464, gl_rom_n_465, gl_rom_n_466, gl_rom_n_467, gl_rom_n_468 : std_logic;
  signal gl_rom_n_469, gl_rom_n_470, gl_rom_n_471, gl_rom_n_472, gl_rom_n_473 : std_logic;
  signal gl_rom_n_474, gl_rom_n_475, gl_rom_n_476, gl_rom_n_477, gl_rom_n_478 : std_logic;
  signal gl_rom_n_479, gl_rom_n_480, gl_rom_n_481, gl_rom_n_482, gl_rom_n_483 : std_logic;
  signal gl_rom_n_484, gl_rom_n_485, gl_rom_n_486, gl_rom_n_487, gl_rom_n_488 : std_logic;
  signal gl_rom_n_489, gl_rom_n_490, gl_rom_n_491, gl_rom_n_492, gl_rom_n_493 : std_logic;
  signal gl_rom_n_494, gl_rom_n_495, gl_rom_n_496, gl_rom_n_497, gl_rom_n_498 : std_logic;
  signal gl_rom_n_499, gl_rom_n_500, gl_rom_n_501, gl_rom_n_502, gl_rom_n_503 : std_logic;
  signal gl_rom_n_504, gl_rom_n_505, gl_rom_n_506, gl_rom_n_507, gl_rom_n_508 : std_logic;
  signal gl_rom_n_509, gl_rom_n_510, gl_rom_n_511, gl_rom_n_512, gl_rom_n_513 : std_logic;
  signal gl_rom_n_514, gl_rom_n_515, gl_rom_n_516, gl_rom_n_517, gl_rom_n_518 : std_logic;
  signal gl_rom_n_519, gl_rom_n_520, gl_rom_n_521, gl_rom_n_522, gl_rom_n_523 : std_logic;
  signal gl_rom_n_524, gl_rom_n_525, gl_rom_n_526, gl_rom_n_527, gl_rom_n_528 : std_logic;
  signal gl_rom_n_529, gl_rom_n_530, gl_rom_n_531, gl_rom_n_532, gl_rom_n_533 : std_logic;
  signal gl_rom_n_534, gl_rom_n_535, gl_rom_n_536, gl_rom_n_537, gl_rom_n_538 : std_logic;
  signal gl_rom_n_539, gl_rom_n_540, gl_rom_n_541, gl_rom_n_542, gl_rom_n_543 : std_logic;
  signal gl_rom_n_544, gl_rom_n_545, gl_rom_n_546, gl_rom_n_547, gl_rom_n_548 : std_logic;
  signal gl_rom_n_549, gl_rom_n_550, gl_rom_n_551, gl_rom_n_552, gl_rom_n_553 : std_logic;
  signal gl_rom_n_554, gl_rom_n_555, gl_rom_n_556, gl_rom_n_557, gl_rom_n_558 : std_logic;
  signal gl_rom_n_559, gl_rom_n_560, gl_rom_n_561, gl_rom_n_562, gl_rom_n_563 : std_logic;
  signal gl_rom_n_564, gl_rom_n_565, gl_rom_n_566, gl_rom_n_567, gl_rom_n_568 : std_logic;
  signal gl_rom_n_569, gl_rom_n_570, gl_rom_n_571, gl_rom_n_572, gl_rom_n_573 : std_logic;
  signal gl_rom_n_574, gl_rom_n_575, gl_rom_n_576, gl_rom_n_577, gl_rom_n_578 : std_logic;
  signal gl_rom_n_579, gl_rom_n_580, gl_rom_n_581, gl_rom_n_582, gl_rom_n_583 : std_logic;
  signal gl_rom_n_584, gl_rom_n_585, gl_rom_n_586, gl_rom_n_587, gl_rom_n_588 : std_logic;
  signal gl_rom_n_589, gl_rom_n_590, gl_rom_n_591, gl_rom_n_592, gl_rom_n_593 : std_logic;
  signal gl_rom_n_594, gl_rom_n_595, gl_rom_n_596, gl_rom_n_597, gl_rom_n_598 : std_logic;
  signal gl_rom_n_599, gl_rom_n_600, gl_rom_n_601, gl_rom_n_602, gl_rom_n_603 : std_logic;
  signal gl_rom_n_604, gl_rom_n_605, gl_rom_n_606, gl_rom_n_607, gl_rom_n_608 : std_logic;
  signal gl_rom_n_609, gl_rom_n_610, gl_rom_n_611, gl_rom_n_612, gl_rom_n_613 : std_logic;
  signal gl_rom_n_614, gl_rom_n_615, gl_rom_n_616, gl_rom_n_617, gl_rom_n_618 : std_logic;
  signal gl_rom_n_619, gl_rom_n_620, gl_rom_n_621, gl_rom_n_622, gl_rom_n_623 : std_logic;
  signal gl_rom_n_624, gl_rom_n_625, gl_rom_n_626, gl_rom_n_627, gl_rom_n_628 : std_logic;
  signal gl_rom_n_629, gl_rom_n_630, gl_rom_n_631, gl_rom_n_632, gl_rom_n_633 : std_logic;
  signal gl_rom_n_634, gl_rom_n_635, gl_rom_n_636, gl_rom_n_637, gl_rom_n_638 : std_logic;
  signal gl_rom_n_639, gl_rom_n_640, gl_rom_n_641, gl_rom_n_642, gl_rom_n_643 : std_logic;
  signal gl_rom_n_644, gl_rom_n_645, gl_rom_n_646, gl_rom_n_647, gl_rom_n_648 : std_logic;
  signal gl_rom_n_649, gl_rom_n_650, gl_rom_n_651, gl_rom_n_652, gl_rom_n_653 : std_logic;
  signal gl_rom_n_654, gl_rom_n_655, gl_rom_n_656, gl_rom_n_657, gl_rom_n_658 : std_logic;
  signal gl_rom_n_659, gl_rom_n_660, gl_rom_n_661, gl_rom_n_662, gl_rom_n_663 : std_logic;
  signal gl_rom_n_664, gl_rom_n_665, gl_rom_n_666, gl_rom_n_667, gl_rom_n_668 : std_logic;
  signal gl_rom_n_669, gl_rom_n_670, gl_rom_n_671, gl_rom_n_672, gl_rom_n_673 : std_logic;
  signal gl_rom_n_674, gl_rom_n_675, gl_rom_n_676, gl_rom_n_677, gl_rom_n_678 : std_logic;
  signal gl_rom_n_679, gl_rom_n_680, gl_rom_n_681, gl_rom_n_682, gl_rom_n_683 : std_logic;
  signal gl_rom_n_684, gl_rom_n_685, gl_rom_n_686, gl_rom_n_687, gl_rom_n_688 : std_logic;
  signal gl_rom_n_689, gl_rom_n_690, gl_rom_n_691, gl_rom_n_692, gl_rom_n_693 : std_logic;
  signal gl_rom_n_694, gl_rom_n_695, gl_rom_n_696, gl_rom_n_697, gl_rom_n_698 : std_logic;
  signal gl_rom_n_699, gl_rom_n_700, gl_rom_n_701, gl_rom_n_702, gl_rom_n_703 : std_logic;
  signal gl_rom_n_704, gl_rom_n_705, gl_rom_n_706, gl_rom_n_707, gl_rom_n_708 : std_logic;
  signal gl_rom_n_709, gl_rom_n_710, gl_rom_n_711, gl_rom_n_712, gl_rom_n_713 : std_logic;
  signal gl_rom_n_714, gl_rom_n_715, gl_rom_n_716, gl_rom_n_717, gl_rom_n_718 : std_logic;
  signal gl_rom_n_719, gl_rom_n_720, gl_rom_n_721, gl_rom_n_722, gl_rom_n_723 : std_logic;
  signal gl_rom_n_724, gl_rom_n_725, gl_rom_n_726, gl_rom_n_727, gl_rom_n_728 : std_logic;
  signal gl_rom_n_729, gl_rom_n_730, gl_rom_n_731, gl_rom_n_732, gl_rom_n_733 : std_logic;
  signal gl_rom_n_734, gl_rom_n_735, gl_rom_n_736, gl_rom_n_737, gl_rom_n_738 : std_logic;
  signal gl_rom_n_739, gl_rom_n_740, gl_rom_n_741, gl_rom_n_742, gl_rom_n_743 : std_logic;
  signal gl_rom_n_744, gl_rom_n_745, gl_rom_n_746, gl_rom_n_747, gl_rom_n_748 : std_logic;
  signal gl_rom_n_749, gl_rom_n_750, gl_rom_n_751, gl_rom_n_752, gl_rom_n_753 : std_logic;
  signal gl_rom_n_754, gl_rom_n_755, gl_rom_n_756, gl_rom_n_757, gl_rom_n_758 : std_logic;
  signal gl_rom_n_759, gl_rom_n_760, gl_rom_n_761, gl_rom_n_762, gl_rom_n_763 : std_logic;
  signal gl_rom_n_764, gl_rom_n_765, gl_rom_n_766, gl_rom_n_767, gl_rom_n_768 : std_logic;
  signal gl_rom_n_769, gl_rom_n_770, gl_rom_n_771, gl_rom_n_772, gl_rom_n_773 : std_logic;
  signal gl_rom_n_774, gl_rom_n_775, gl_rom_n_776, gl_rom_n_777, gl_rom_n_778 : std_logic;
  signal gl_rom_n_779, gl_rom_n_780, gl_rom_n_781, gl_rom_n_782, gl_rom_n_783 : std_logic;
  signal gl_rom_n_784, gl_rom_n_785, gl_rom_n_786, gl_rom_n_787, gl_rom_n_788 : std_logic;
  signal gl_rom_n_789, gl_rom_n_790, gl_rom_n_791, gl_rom_n_792, gl_rom_n_793 : std_logic;
  signal gl_rom_n_794, gl_rom_n_795, gl_rom_n_796, gl_rom_n_797, gl_rom_n_798 : std_logic;
  signal gl_rom_n_799, gl_rom_n_800, gl_rom_n_801, gl_rom_n_802, gl_rom_n_803 : std_logic;
  signal gl_rom_n_804, gl_rom_n_805, gl_rom_n_806, gl_rom_n_807, gl_rom_n_808 : std_logic;
  signal gl_rom_n_809, gl_rom_n_810, gl_rom_n_811, gl_rom_n_812, gl_rom_n_813 : std_logic;
  signal gl_rom_n_814, gl_rom_n_815, gl_rom_n_816, gl_rom_n_817, gl_rom_n_818 : std_logic;
  signal gl_rom_n_819, gl_rom_n_820, gl_rom_n_821, gl_rom_n_822, gl_rom_n_823 : std_logic;
  signal gl_rom_n_824, gl_rom_n_825, gl_rom_n_826, gl_rom_n_827, gl_rom_n_828 : std_logic;
  signal gl_rom_n_829, gl_rom_n_830, gl_rom_n_831, gl_rom_n_832, gl_rom_n_833 : std_logic;
  signal gl_rom_n_834, gl_rom_n_835, gl_rom_n_836, gl_rom_n_837, gl_rom_n_838 : std_logic;
  signal gl_rom_n_839, gl_rom_n_840, gl_rom_n_841, gl_rom_n_842, gl_rom_n_843 : std_logic;
  signal gl_rom_n_844, gl_rom_n_845, gl_rom_n_846, gl_rom_n_847, gl_rom_n_848 : std_logic;
  signal gl_rom_n_849, gl_rom_n_850, gl_rom_n_851, gl_rom_n_852, gl_rom_n_853 : std_logic;
  signal gl_rom_n_854, gl_rom_n_855, gl_rom_n_856, gl_rom_n_857, gl_rom_n_858 : std_logic;
  signal gl_rom_n_859, gl_rom_n_860, gl_rom_n_861, gl_rom_n_862, gl_rom_n_863 : std_logic;
  signal gl_rom_n_864, gl_rom_n_865, gl_rom_n_866, gl_rom_n_867, gl_rom_n_868 : std_logic;
  signal gl_rom_n_869, gl_rom_n_870, gl_rom_n_871, gl_rom_n_872, gl_rom_n_873 : std_logic;
  signal gl_rom_n_874, gl_rom_n_875, gl_rom_n_876, gl_rom_n_877, gl_rom_n_878 : std_logic;
  signal gl_rom_n_879, gl_rom_n_880, gl_rom_n_881, gl_rom_n_882, gl_rom_n_883 : std_logic;
  signal gl_rom_n_884, gl_rom_n_885, gl_rom_n_886, gl_rom_n_887, gl_rom_n_888 : std_logic;
  signal gl_rom_n_889, gl_rom_n_890, gl_rom_n_891, gl_rom_n_892, gl_rom_n_893 : std_logic;
  signal gl_rom_n_894, gl_rom_n_895, gl_rom_n_896, gl_rom_n_897, gl_rom_n_898 : std_logic;
  signal gl_rom_n_899, gl_rom_n_900, gl_rom_n_901, gl_rom_n_902, gl_rom_n_903 : std_logic;
  signal gl_rom_n_904, gl_rom_n_905, gl_rom_n_906, gl_rom_n_907, gl_rom_n_908 : std_logic;
  signal gl_rom_n_909, gl_rom_n_910, gl_rom_n_911, gl_rom_n_912, gl_rom_n_913 : std_logic;
  signal gl_rom_n_914, gl_rom_n_915, gl_rom_n_916, gl_rom_n_917, gl_rom_n_918 : std_logic;
  signal gl_rom_n_919, gl_rom_n_920, gl_rom_n_921, gl_rom_n_922, gl_rom_n_923 : std_logic;
  signal gl_rom_n_924, gl_rom_n_925, gl_rom_n_926, gl_rom_n_927, gl_rom_n_928 : std_logic;
  signal gl_rom_n_929, gl_rom_n_930, gl_rom_n_931, gl_rom_n_932, gl_rom_n_933 : std_logic;
  signal gl_rom_n_934, gl_rom_n_935, gl_rom_n_936, gl_rom_n_937, gl_rom_n_938 : std_logic;
  signal gl_rom_n_939, gl_rom_n_940, gl_rom_n_941, gl_rom_n_942, gl_rom_n_943 : std_logic;
  signal gl_rom_n_944, gl_rom_n_945, gl_rom_n_946, gl_rom_n_947, gl_rom_n_948 : std_logic;
  signal gl_rom_n_949, gl_rom_n_950, gl_rom_n_951, gl_rom_n_952, gl_rom_n_953 : std_logic;
  signal gl_rom_n_954, gl_rom_n_955, gl_rom_n_956, gl_rom_n_957, gl_rom_n_958 : std_logic;
  signal gl_rom_n_959, gl_rom_n_960, gl_rom_n_961, gl_rom_n_962, gl_rom_n_963 : std_logic;
  signal gl_rom_n_964, gl_rom_n_965, gl_rom_n_966, gl_rom_n_967, gl_rom_n_968 : std_logic;
  signal gl_rom_n_969, gl_rom_n_970, gl_rom_n_971, gl_rom_n_972, gl_rom_n_973 : std_logic;
  signal gl_rom_n_974, gl_rom_n_975, gl_rom_n_976, gl_rom_n_977, gl_rom_n_978 : std_logic;
  signal gl_rom_n_979, gl_rom_n_980, gl_rom_n_981, gl_rom_n_982, gl_rom_n_983 : std_logic;
  signal gl_rom_n_984, gl_rom_n_985, gl_rom_n_986, gl_rom_n_987, gl_rom_n_988 : std_logic;
  signal gl_rom_n_989, gl_rom_n_990, gl_rom_n_991, gl_rom_n_992, gl_rom_n_993 : std_logic;
  signal gl_rom_n_994, gl_rom_n_995, gl_rom_n_996, gl_rom_n_997, gl_rom_n_998 : std_logic;
  signal gl_rom_n_999, gl_rom_n_1000, gl_rom_n_1001, gl_rom_n_1002, gl_rom_n_1003 : std_logic;
  signal gl_rom_n_1004, gl_rom_n_1005, gl_rom_n_1006, gl_rom_n_1007, gl_rom_n_1008 : std_logic;
  signal gl_rom_n_1009, gl_rom_n_1010, gl_rom_n_1011, gl_rom_n_1012, gl_rom_n_1013 : std_logic;
  signal gl_rom_n_1014, gl_rom_n_1015, gl_rom_n_1016, gl_rom_n_1017, gl_rom_n_1018 : std_logic;
  signal gl_rom_n_1019, gl_rom_n_1020, gl_rom_n_1021, gl_rom_n_1022, gl_rom_n_1023 : std_logic;
  signal gl_rom_n_1024, gl_rom_n_1025, gl_rom_n_1026, gl_rom_n_1027, gl_rom_n_1028 : std_logic;
  signal gl_rom_n_1029, gl_rom_n_1030, gl_rom_n_1031, gl_rom_n_1032, gl_rom_n_1033 : std_logic;
  signal gl_rom_n_1034, gl_rom_n_1035, gl_rom_n_1036, gl_rom_n_1037, gl_rom_n_1038 : std_logic;
  signal gl_rom_n_1039, gl_rom_n_1040, gl_rom_n_1041, gl_rom_n_1042, gl_rom_n_1043 : std_logic;
  signal gl_rom_n_1044, gl_rom_n_1045, gl_rom_n_1046, gl_rom_n_1047, gl_rom_n_1048 : std_logic;
  signal gl_rom_n_1049, gl_rom_n_1050, gl_rom_n_1051, gl_rom_n_1052, gl_rom_n_1053 : std_logic;
  signal gl_rom_n_1054, gl_rom_n_1055, gl_rom_n_1056, gl_rom_n_1057, gl_rom_n_1058 : std_logic;
  signal gl_rom_n_1059, gl_rom_n_1060, gl_rom_n_1061, gl_rom_n_1062, gl_rom_n_1063 : std_logic;
  signal gl_rom_n_1064, gl_rom_n_1065, gl_rom_n_1066, gl_rom_n_1067, gl_rom_n_1068 : std_logic;
  signal gl_rom_n_1069, gl_rom_n_1070, gl_rom_n_1071, gl_rom_n_1072, gl_rom_n_1073 : std_logic;
  signal gl_rom_n_1074, gl_rom_n_1075, gl_rom_n_1076, gl_rom_n_1077, gl_rom_n_1078 : std_logic;
  signal gl_rom_n_1079, gl_rom_n_1080, gl_rom_n_1081, gl_rom_n_1082, gl_rom_n_1083 : std_logic;
  signal gl_rom_n_1084, gl_rom_n_1085, gl_rom_n_1086, gl_rom_n_1087, gl_rom_n_1088 : std_logic;
  signal gl_rom_n_1089, gl_rom_n_1090, gl_rom_n_1091, gl_rom_n_1092, gl_rom_n_1093 : std_logic;
  signal gl_rom_n_1094, gl_rom_n_1095, gl_rom_n_1096, gl_rom_n_1097, gl_rom_n_1098 : std_logic;
  signal gl_rom_n_1099, gl_rom_n_1100, gl_rom_n_1101, gl_rom_n_1102, gl_rom_n_1103 : std_logic;
  signal gl_rom_n_1104, gl_rom_n_1105, gl_rom_n_1106, gl_rom_n_1107, gl_rom_n_1108 : std_logic;
  signal gl_rom_n_1109, gl_rom_n_1110, gl_rom_n_1111, gl_rom_n_1112, gl_rom_n_1113 : std_logic;
  signal gl_rom_n_1114, gl_rom_n_1115, gl_rom_n_1116, gl_rom_n_1117, gl_rom_n_1118 : std_logic;
  signal gl_rom_n_1119, gl_rom_n_1120, gl_rom_n_1121, gl_rom_n_1122, gl_rom_n_1123 : std_logic;
  signal gl_rom_n_1124, gl_rom_n_1125, gl_rom_n_1126, gl_rom_n_1127, gl_rom_n_1128 : std_logic;
  signal gl_rom_n_1129, gl_rom_n_1130, gl_rom_n_1131, gl_rom_n_1132, gl_rom_n_1133 : std_logic;
  signal gl_rom_n_1134, gl_rom_n_1135, gl_rom_n_1136, gl_rom_n_1137, gl_rom_n_1138 : std_logic;
  signal gl_rom_n_1139, gl_rom_n_1140, gl_rom_n_1141, gl_rom_n_1142, gl_rom_n_1143 : std_logic;
  signal gl_rom_n_1144, gl_rom_n_1145, gl_rom_n_1146, gl_rom_n_1147, gl_rom_n_1148 : std_logic;
  signal gl_rom_n_1149, gl_rom_n_1150, gl_rom_n_1151, gl_rom_n_1152, gl_rom_n_1153 : std_logic;
  signal gl_rom_n_1154, gl_rom_n_1155, gl_rom_n_1156, gl_rom_n_1157, gl_rom_n_1158 : std_logic;
  signal gl_rom_n_1159, gl_rom_n_1160, gl_rom_n_1161, gl_rom_n_1162, gl_rom_n_1163 : std_logic;
  signal gl_rom_n_1164, gl_rom_n_1165, gl_rom_n_1166, gl_rom_n_1167, gl_rom_n_1168 : std_logic;
  signal gl_rom_n_1169, gl_rom_n_1170, gl_rom_n_1171, gl_rom_n_1172, gl_rom_n_1173 : std_logic;
  signal gl_rom_n_1174, gl_rom_n_1175, gl_rom_n_1176, gl_rom_n_1177, gl_rom_n_1178 : std_logic;
  signal gl_rom_n_1179, gl_rom_n_1180, gl_rom_n_1181, gl_rom_n_1182, gl_rom_n_1183 : std_logic;
  signal gl_rom_n_1184, gl_rom_n_1185, gl_rom_n_1186, gl_rom_n_1187, gl_rom_n_1188 : std_logic;
  signal gl_rom_n_1189, gl_rom_n_1190, gl_rom_n_1191, gl_rom_n_1192, gl_rom_n_1193 : std_logic;
  signal gl_rom_n_1194, gl_rom_n_1195, gl_rom_n_1196, gl_rom_n_1197, gl_rom_n_1198 : std_logic;
  signal gl_rom_n_1199, gl_rom_n_1200, gl_rom_n_1201, gl_rom_n_1202, gl_rom_n_1203 : std_logic;
  signal gl_rom_n_1204, gl_rom_n_1205, gl_rom_n_1206, gl_rom_n_1207, gl_rom_n_1208 : std_logic;
  signal gl_rom_n_1209, gl_rom_n_1210, gl_rom_n_1211, gl_rom_n_1212, gl_rom_n_1213 : std_logic;
  signal gl_rom_n_1214, gl_rom_n_1215, gl_rom_n_1216, gl_rom_n_1217, gl_rom_n_1218 : std_logic;
  signal gl_rom_n_1219, gl_rom_n_1220, gl_rom_n_1221, gl_rom_n_1222, gl_rom_n_1223 : std_logic;
  signal gl_rom_n_1224, gl_rom_n_1225, gl_rom_n_1226, gl_rom_n_1227, gl_rom_n_1228 : std_logic;
  signal gl_rom_n_1229, gl_rom_n_1230, gl_rom_n_1231, gl_rom_n_1232, gl_rom_n_1233 : std_logic;
  signal gl_rom_n_1234, gl_rom_n_1235, gl_rom_n_1236, gl_rom_n_1237, gl_rom_n_1238 : std_logic;
  signal gl_rom_n_1239, gl_rom_n_1240, gl_rom_n_1241, gl_rom_n_1242, gl_rom_n_1243 : std_logic;
  signal gl_rom_n_1244, gl_rom_n_1245, gl_rom_n_1246, gl_rom_n_1247, gl_rom_n_1248 : std_logic;
  signal gl_rom_n_1249, gl_rom_n_1250, gl_rom_n_1251, gl_rom_n_1252, gl_rom_n_1253 : std_logic;
  signal gl_rom_n_1254, gl_rom_n_1255, gl_rom_n_1256, gl_rom_n_1257, gl_rom_n_1258 : std_logic;
  signal gl_rom_n_1259, gl_rom_n_1260, gl_rom_n_1261, gl_rom_n_1262, gl_rom_n_1263 : std_logic;
  signal gl_rom_n_1264, gl_rom_n_1265, gl_rom_n_1266, gl_rom_n_1267, gl_rom_n_1268 : std_logic;
  signal gl_rom_n_1269, gl_rom_n_1270, gl_rom_n_1271, gl_rom_n_1272, gl_rom_n_1273 : std_logic;
  signal gl_rom_n_1274, gl_rom_n_1275, gl_rom_n_1276, gl_rom_n_1277, gl_rom_n_1278 : std_logic;
  signal gl_rom_n_1279, gl_rom_n_1280, gl_rom_n_1281, gl_rom_n_1282, gl_rom_n_1283 : std_logic;
  signal gl_rom_n_1284, gl_rom_n_1285, gl_rom_n_1286, gl_rom_n_1287, gl_rom_n_1288 : std_logic;
  signal gl_rom_n_1289, gl_rom_n_1290, gl_rom_n_1291, gl_rom_n_1292, gl_rom_n_1293 : std_logic;
  signal gl_rom_n_1294, gl_rom_n_1295, gl_rom_n_1296, gl_rom_n_1297, gl_rom_n_1298 : std_logic;
  signal gl_rom_n_1299, gl_rom_n_1300, gl_rom_n_1301, gl_rom_n_1302, gl_rom_n_1303 : std_logic;
  signal gl_rom_n_1304, gl_rom_n_1305, gl_rom_n_1306, gl_rom_n_1307, gl_rom_n_1308 : std_logic;
  signal gl_rom_n_1309, gl_rom_n_1310, gl_rom_n_1311, gl_rom_n_1312, gl_rom_n_1313 : std_logic;
  signal gl_rom_n_1314, gl_rom_n_1315, gl_rom_n_1316, gl_rom_n_1317, gl_rom_n_1318 : std_logic;
  signal gl_rom_n_1319, gl_rom_n_1320, gl_rom_n_1321, gl_rom_n_1322, gl_rom_n_1323 : std_logic;
  signal gl_rom_n_1324, gl_rom_n_1325, gl_rom_n_1326, gl_rom_n_1327, gl_rom_n_1328 : std_logic;
  signal gl_rom_n_1329, gl_rom_n_1330, gl_rom_n_1331, gl_rom_n_1332, gl_rom_n_1333 : std_logic;
  signal gl_rom_n_1334, gl_rom_n_1335, gl_rom_n_1336, gl_rom_n_1337, gl_rom_n_1338 : std_logic;
  signal gl_rom_n_1339, gl_rom_n_1340, gl_rom_n_1341, gl_rom_n_1342, gl_rom_n_1343 : std_logic;
  signal gl_rom_n_1344, gl_rom_n_1345, gl_rom_n_1346, gl_rom_n_1347, gl_rom_n_1348 : std_logic;
  signal gl_rom_n_1349, gl_rom_n_1350, gl_rom_n_1351, gl_rom_n_1352, gl_rom_n_1353 : std_logic;
  signal gl_rom_n_1354, gl_rom_n_1355, gl_rom_n_1356, gl_rom_n_1357, gl_rom_n_1358 : std_logic;
  signal gl_rom_n_1359, gl_rom_n_1360, gl_rom_n_1361, gl_rom_n_1362, gl_rom_n_1363 : std_logic;
  signal gl_rom_n_1364, gl_rom_n_1365, gl_rom_n_1366, gl_rom_n_1367, gl_rom_n_1368 : std_logic;
  signal gl_rom_n_1369, gl_rom_n_1370, gl_rom_n_1371, gl_rom_n_1372, gl_rom_n_1373 : std_logic;
  signal gl_rom_n_1374, gl_rom_n_1375, gl_rom_n_1376, gl_rom_n_1377, gl_rom_n_1378 : std_logic;
  signal gl_rom_n_1379, gl_rom_n_1380, gl_rom_n_1381, gl_rom_n_1382, gl_rom_n_1383 : std_logic;
  signal gl_rom_n_1384, gl_rom_n_1385, gl_rom_n_1386, gl_rom_n_1387, gl_rom_n_1388 : std_logic;
  signal gl_rom_n_1389, gl_rom_n_1390, gl_rom_n_1391, gl_rom_n_1392, gl_rom_n_1393 : std_logic;
  signal gl_rom_n_1394, gl_rom_n_1395, gl_rom_n_1396, gl_rom_n_1397, gl_rom_n_1398 : std_logic;
  signal gl_rom_n_1399, gl_rom_n_1400, gl_rom_n_1401, gl_rom_n_1402, gl_rom_n_1403 : std_logic;
  signal gl_rom_n_1404, gl_rom_n_1405, gl_rom_n_1406, gl_rom_n_1407, gl_rom_n_1408 : std_logic;
  signal gl_rom_n_1409, gl_rom_n_1410, gl_rom_n_1411, gl_rom_n_1412, gl_rom_n_1413 : std_logic;
  signal gl_rom_n_1414, gl_rom_n_1415, gl_rom_n_1416, gl_rom_n_1417, gl_rom_n_1418 : std_logic;
  signal gl_rom_n_1419, gl_rom_n_1420, gl_rom_n_1421, gl_rom_n_1422, gl_rom_n_1423 : std_logic;
  signal gl_rom_n_1424, gl_rom_n_1425, gl_rom_n_1426, gl_rom_n_1427, gl_rom_n_1428 : std_logic;
  signal gl_rom_n_1429, gl_rom_n_1430, gl_rom_n_1431, gl_rom_n_1432, gl_rom_n_1433 : std_logic;
  signal gl_rom_n_1434, gl_rom_n_1435, gl_rom_n_1436, gl_rom_n_1437, gl_rom_n_1438 : std_logic;
  signal gl_rom_n_1439, gl_rom_n_1440, gl_rom_n_1441, gl_rom_n_1442, gl_rom_n_1443 : std_logic;
  signal gl_rom_n_1444, gl_rom_n_1445, gl_rom_n_1446, gl_rom_n_1447, gl_rom_n_1448 : std_logic;
  signal gl_rom_n_1449, gl_rom_n_1450, gl_rom_n_1451, gl_rom_n_1452, gl_rom_n_1453 : std_logic;
  signal gl_rom_n_1454, gl_rom_n_1455, gl_rom_n_1456, gl_rom_n_1457, gl_rom_n_1458 : std_logic;
  signal gl_rom_n_1459, gl_rom_n_1460, gl_rom_n_1461, gl_rom_n_1462, gl_rom_n_1463 : std_logic;
  signal gl_rom_n_1464, gl_rom_n_1465, gl_rom_n_1466, gl_rom_n_1467, gl_rom_n_1468 : std_logic;
  signal gl_rom_n_1469, gl_rom_n_1470, gl_rom_n_1471, gl_rom_n_1472, gl_rom_n_1473 : std_logic;
  signal gl_rom_n_1474, gl_rom_n_1475, gl_rom_n_1476, gl_rom_n_1477, gl_rom_n_1478 : std_logic;
  signal gl_rom_n_1479, gl_rom_n_1480, gl_rom_n_1481, gl_rom_n_1482, gl_rom_n_1483 : std_logic;
  signal gl_rom_n_1484, gl_rom_n_1485, gl_rom_n_1486, gl_rom_n_1487, gl_rom_n_1488 : std_logic;
  signal gl_rom_n_1489, gl_rom_n_1490, gl_rom_n_1491, gl_rom_n_1492, gl_rom_n_1493 : std_logic;
  signal gl_rom_n_1494, gl_rom_n_1495, gl_rom_n_1496, gl_rom_n_1497, gl_rom_n_1498 : std_logic;
  signal gl_rom_n_1499, gl_rom_n_1500, gl_sig_blue, gl_sig_green, gl_sig_red : std_logic;
  signal gl_sig_scale_h, gl_sig_scale_v, gl_vgd_n_0, gl_vgd_n_2, gl_vgd_n_3 : std_logic;
  signal gl_vgd_n_4, gl_vgd_n_5, gl_vgd_n_6, gl_vgd_n_7, gl_vgd_n_8 : std_logic;
  signal gl_vgd_n_9, gl_vgd_n_10, gl_vgd_n_11, gl_vgd_n_12, gl_vgd_n_13 : std_logic;
  signal gl_vgd_n_14, gl_vgd_n_15, gl_vgd_n_16, gl_vgd_n_17, gl_vgd_n_18 : std_logic;
  signal gl_vgd_n_19, gl_vgd_n_20, gl_vgd_n_21, gl_vgd_n_22, gl_vgd_n_23 : std_logic;
  signal gl_vgd_n_24, gl_vgd_n_25, gl_vgd_n_26, gl_vgd_n_27, gl_vgd_n_28 : std_logic;
  signal gl_vgd_n_29, gl_vgd_n_30, gl_vgd_n_31, gl_vgd_n_32, gl_vgd_n_33 : std_logic;
  signal gl_vgd_n_34, gl_vgd_n_35, gl_vgd_n_36, gl_vgd_n_37, gl_vgd_n_38 : std_logic;
  signal gl_vgd_n_39, gl_vgd_n_40, gl_vgd_n_41, gl_vgd_n_42, gl_vgd_n_43 : std_logic;
  signal gl_vgd_n_44, gl_vgd_n_45, gl_vgd_n_46, gl_vgd_n_47, gl_vgd_n_48 : std_logic;
  signal gl_vgd_n_49, gl_vgd_n_50, gl_vgd_n_51, gl_vgd_n_52, gl_vgd_n_53 : std_logic;
  signal gl_vgd_n_54, gl_vgd_n_55, gl_vgd_n_56, gl_vgd_n_57, gl_vgd_n_58 : std_logic;
  signal gl_vgd_n_59, gl_vgd_n_60, gl_vgd_n_61, gl_vgd_n_62, gl_vgd_n_63 : std_logic;
  signal gl_vgd_n_64, gl_vgd_n_65, gl_vgd_n_67, gl_vgd_n_68, gl_vgd_n_69 : std_logic;
  signal gl_vgd_n_70, gl_vgd_n_71, gl_vgd_n_72, gl_vgd_n_73, gl_vgd_n_74 : std_logic;
  signal gl_vgd_n_75, gl_vgd_n_76, gl_vgd_n_77, gl_vgd_n_78, gl_vgd_n_79 : std_logic;
  signal gl_vgd_n_80, gl_vgd_n_81, gl_vgd_n_82, gl_vgd_n_83, logic_1_1_net : std_logic;
  signal ml_handshake_mouse_out, ml_il_color1_n_0, ml_il_color1_n_1, ml_il_color1_n_3, ml_il_color1_n_4 : std_logic;
  signal ml_il_color1_n_5, ml_il_color1_n_6, ml_il_color1_n_7, ml_il_color1_n_8, ml_il_color1_n_9 : std_logic;
  signal ml_il_color1_n_10, ml_il_color1_n_11, ml_il_color1_n_12, ml_il_color1_n_14, ml_il_color1_n_15 : std_logic;
  signal ml_il_color1_n_16, ml_il_color1_n_17, ml_il_color1_n_18, ml_il_color1_n_20, ml_il_color1_n_21 : std_logic;
  signal ml_il_color1_n_22, ml_il_color1_n_23, ml_il_x1_n_1, ml_il_x1_n_2, ml_il_x1_n_3 : std_logic;
  signal ml_il_x1_n_4, ml_il_x1_n_5, ml_il_x1_n_6, ml_il_x1_n_7, ml_il_x1_n_8 : std_logic;
  signal ml_il_x1_n_9, ml_il_x1_n_13, ml_il_x1_n_14, ml_il_x1_n_15, ml_il_x1_n_16 : std_logic;
  signal ml_il_x1_n_17, ml_il_x1_n_18, ml_il_x1_n_19, ml_il_x1_n_20, ml_il_x1_n_21 : std_logic;
  signal ml_il_x1_n_22, ml_il_x1_n_23, ml_il_x1_n_24, ml_il_x1_n_25, ml_il_x1_n_26 : std_logic;
  signal ml_il_x1_n_27, ml_il_x1_n_28, ml_il_x1_n_29, ml_il_x1_n_39, ml_il_x1_n_40 : std_logic;
  signal ml_il_x1_n_41, ml_il_x1_n_42, ml_il_x1_n_43, ml_il_x1_n_47, ml_il_x1_n_48 : std_logic;
  signal ml_il_x1_n_49, ml_il_y1_n_1, ml_il_y1_n_2, ml_il_y1_n_3, ml_il_y1_n_4 : std_logic;
  signal ml_il_y1_n_5, ml_il_y1_n_6, ml_il_y1_n_7, ml_il_y1_n_8, ml_il_y1_n_9 : std_logic;
  signal ml_il_y1_n_13, ml_il_y1_n_14, ml_il_y1_n_15, ml_il_y1_n_16, ml_il_y1_n_17 : std_logic;
  signal ml_il_y1_n_18, ml_il_y1_n_19, ml_il_y1_n_20, ml_il_y1_n_21, ml_il_y1_n_22 : std_logic;
  signal ml_il_y1_n_23, ml_il_y1_n_24, ml_il_y1_n_25, ml_il_y1_n_26, ml_il_y1_n_27 : std_logic;
  signal ml_il_y1_n_28, ml_il_y1_n_29, ml_il_y1_n_39, ml_il_y1_n_40, ml_il_y1_n_41 : std_logic;
  signal ml_il_y1_n_42, ml_il_y1_n_43, ml_il_y1_n_47, ml_il_y1_n_48, ml_il_y1_n_49 : std_logic;
  signal ml_ms_actBit, ml_ms_btnflipfloprst, ml_ms_cntD_n_0, ml_ms_cntD_n_1, ml_ms_cntD_n_2 : std_logic;
  signal ml_ms_cntD_n_3, ml_ms_cntD_n_4, ml_ms_cntD_n_5, ml_ms_cntD_n_6, ml_ms_cntD_n_7 : std_logic;
  signal ml_ms_cntD_n_8, ml_ms_cntD_n_9, ml_ms_cntD_n_10, ml_ms_cntD_n_11, ml_ms_cntD_n_12 : std_logic;
  signal ml_ms_cntD_n_13, ml_ms_cntD_n_14, ml_ms_cntD_n_15, ml_ms_cntD_n_16, ml_ms_cntD_n_17 : std_logic;
  signal ml_ms_cntD_n_18, ml_ms_cntD_n_19, ml_ms_cntD_n_20, ml_ms_cntD_n_21, ml_ms_cntD_n_22 : std_logic;
  signal ml_ms_cntD_n_23, ml_ms_cntReset15K, ml_ms_cntReset25M, ml_ms_cntReset25M_main, ml_ms_cntReset25M_send : std_logic;
  signal ml_ms_cnt_n_0, ml_ms_cnt_n_1, ml_ms_cnt_n_2, ml_ms_cnt_n_3, ml_ms_cnt_n_4 : std_logic;
  signal ml_ms_cnt_n_5, ml_ms_cnt_n_6, ml_ms_cnt_n_7, ml_ms_cnt_n_8, ml_ms_cnt_n_9 : std_logic;
  signal ml_ms_cnt_n_10, ml_ms_cnt_n_11, ml_ms_cnt_n_12, ml_ms_cnt_n_13, ml_ms_cnt_n_14 : std_logic;
  signal ml_ms_cnt_n_15, ml_ms_cnt_n_16, ml_ms_cnt_n_17, ml_ms_cnt_n_18, ml_ms_cnt_n_19 : std_logic;
  signal ml_ms_cnt_n_20, ml_ms_cnt_n_21, ml_ms_cnt_n_22, ml_ms_cnt_n_23, ml_ms_count_debounce_reset : std_logic;
  signal ml_ms_ed_n_0, ml_ms_ed_n_1, ml_ms_ed_n_2, ml_ms_ed_n_3, ml_ms_ed_n_4 : std_logic;
  signal ml_ms_ed_n_5, ml_ms_ed_n_6, ml_ms_ed_n_7, ml_ms_ed_n_8, ml_ms_ed_n_9 : std_logic;
  signal ml_ms_ed_reg1, ml_ms_ed_reg2, ml_ms_mfsm_n_0, ml_ms_mfsm_n_1, ml_ms_mfsm_n_2 : std_logic;
  signal ml_ms_mfsm_n_4, ml_ms_mfsm_n_5, ml_ms_mfsm_n_6, ml_ms_mfsm_n_7, ml_ms_mfsm_n_8 : std_logic;
  signal ml_ms_mfsm_n_9, ml_ms_mfsm_n_10, ml_ms_mfsm_n_11, ml_ms_mfsm_n_12, ml_ms_mfsm_n_14 : std_logic;
  signal ml_ms_mfsm_n_15, ml_ms_mfsm_n_16, ml_ms_mfsm_n_17, ml_ms_mfsm_n_18, ml_ms_mfsm_n_19 : std_logic;
  signal ml_ms_mfsm_n_20, ml_ms_mfsm_n_21, ml_ms_mfsm_n_22, ml_ms_mfsm_n_23, ml_ms_mfsm_n_24 : std_logic;
  signal ml_ms_mfsm_n_25, ml_ms_mfsm_n_26, ml_ms_mfsm_n_27, ml_ms_mfsm_n_28, ml_ms_mfsm_n_29 : std_logic;
  signal ml_ms_mfsm_n_30, ml_ms_mfsm_n_31, ml_ms_mfsm_n_32, ml_ms_mfsm_n_33, ml_ms_mfsm_n_34 : std_logic;
  signal ml_ms_mfsm_n_35, ml_ms_mfsm_n_36, ml_ms_mfsm_n_37, ml_ms_mfsm_n_38, ml_ms_mfsm_n_39 : std_logic;
  signal ml_ms_mfsm_n_40, ml_ms_mfsm_n_41, ml_ms_mfsm_n_42, ml_ms_mfsm_n_43, ml_ms_mfsm_n_44 : std_logic;
  signal ml_ms_mfsm_n_45, ml_ms_mfsm_n_46, ml_ms_mfsm_n_47, ml_ms_mfsm_n_48, ml_ms_mfsm_n_49 : std_logic;
  signal ml_ms_mfsm_n_50, ml_ms_mfsm_n_51, ml_ms_mfsm_n_52, ml_ms_mfsm_n_53, ml_ms_mfsm_n_54 : std_logic;
  signal ml_ms_mfsm_n_55, ml_ms_mfsm_n_56, ml_ms_mfsm_n_57, ml_ms_mfsm_n_57_BAR, ml_ms_mfsm_n_58 : std_logic;
  signal ml_ms_mfsm_n_60, ml_ms_mfsm_n_108, ml_ms_mfsm_n_109, ml_ms_mfsm_n_110, ml_ms_muxFSM : std_logic;
  signal ml_ms_muxReg, ml_ms_mux_select, ml_ms_mux_select_main, ml_ms_mx_n_0, ml_ms_mx_n_1 : std_logic;
  signal ml_ms_n_0, ml_ms_n_1, ml_ms_n_2, ml_ms_n_3, ml_ms_n_4 : std_logic;
  signal ml_ms_n_5, ml_ms_n_6, ml_ms_n_7, ml_ms_n_8, ml_ms_n_9 : std_logic;
  signal ml_ms_n_10, ml_ms_n_11, ml_ms_n_12, ml_ms_n_13, ml_ms_n_14 : std_logic;
  signal ml_ms_n_15, ml_ms_n_16, ml_ms_n_17, ml_ms_n_18, ml_ms_n_19 : std_logic;
  signal ml_ms_n_20, ml_ms_n_21, ml_ms_n_22, ml_ms_n_23, ml_ms_n_24 : std_logic;
  signal ml_ms_n_25, ml_ms_n_26, ml_ms_n_27, ml_ms_n_28, ml_ms_n_29 : std_logic;
  signal ml_ms_n_30, ml_ms_n_31, ml_ms_n_32, ml_ms_n_33, ml_ms_n_34 : std_logic;
  signal ml_ms_n_35, ml_ms_n_36, ml_ms_n_37, ml_ms_n_38, ml_ms_n_39 : std_logic;
  signal ml_ms_n_40, ml_ms_n_41, ml_ms_n_42, ml_ms_n_43, ml_ms_n_44 : std_logic;
  signal ml_ms_n_45, ml_ms_n_46, ml_ms_n_47, ml_ms_n_48, ml_ms_n_49 : std_logic;
  signal ml_ms_n_50, ml_ms_n_51, ml_ms_n_52, ml_ms_n_53, ml_ms_n_54 : std_logic;
  signal ml_ms_n_55, ml_ms_n_56, ml_ms_n_57, ml_ms_n_58, ml_ms_n_59 : std_logic;
  signal ml_ms_n_60, ml_ms_n_61, ml_ms_n_62, ml_ms_n_63, ml_ms_output_edgedet : std_logic;
  signal ml_ms_reset_send, ml_ms_sfsm_n_383, ml_ms_sr11_data_out_0_79, ml_ms_sr11_data_out_1_80, ml_ms_sr11_data_out_5_84 : std_logic;
  signal ml_ms_tb_n_0, ml_ms_tb_n_1, ml_ms_tb_n_2, ml_ms_tb_n_3, ml_ms_tb_n_4 : std_logic;
  signal ml_ms_tb_n_5, ml_ms_tb_n_6, ml_ms_xflipfloprst, ml_ms_yflipfloprst, sig_countlow : std_logic;
  signal sig_draw, sig_rescount : std_logic;

begin

  FE_PHC530_sig_logic_y_2 : BUFFD1BWP7T port map(I => FE_PHN525_sig_logic_y_2, Z => FE_PHN530_sig_logic_y_2);
  FE_PHC529_sig_logic_y_1 : DEL01BWP7T port map(I => sig_logic_y(1), Z => FE_PHN529_sig_logic_y_1);
  FE_PHC528_sig_logic_y_3 : CKBD1BWP7T port map(I => FE_PHN316_sig_logic_y_3, Z => FE_PHN528_sig_logic_y_3);
  FE_PHC527_sig_logic_x_3 : CKBD1BWP7T port map(I => FE_PHN524_sig_logic_x_3, Z => FE_PHN527_sig_logic_x_3);
  FE_PHC526_gl_ram_n_819 : CKBD1BWP7T port map(I => FE_PHN285_gl_ram_n_819, Z => FE_PHN526_gl_ram_n_819);
  FE_PHC525_sig_logic_y_2 : DEL015BWP7T port map(I => sig_logic_y(2), Z => FE_PHN525_sig_logic_y_2);
  FE_PHC524_sig_logic_x_3 : CKBD0BWP7T port map(I => FE_PHN287_sig_logic_x_3, Z => FE_PHN524_sig_logic_x_3);
  FE_PHC523_sig_logic_y_3 : BUFFD0BWP7T port map(I => FE_PHN528_sig_logic_y_3, Z => FE_PHN523_sig_logic_y_3);
  FE_PHC522_FE_OFN4_gl_ram_n_1111 : CKBD8BWP7T port map(I => FE_PHN326_FE_OFN4_gl_ram_n_1111, Z => FE_PHN522_FE_OFN4_gl_ram_n_1111);
  FE_PHC521_gl_ram_n_1111 : BUFFD1P5BWP7T port map(I => FE_PHN521_gl_ram_n_1111, Z => FE_PHN301_gl_ram_n_1111);
  FE_PHC520_gl_ram_n_1111 : DEL01BWP7T port map(I => FE_PHN302_gl_ram_n_1111, Z => FE_PHN520_gl_ram_n_1111);
  FE_PHC519_gl_ram_n_819 : CKBD0BWP7T port map(I => FE_PHN526_gl_ram_n_819, Z => FE_PHN519_gl_ram_n_819);
  FE_PHC518_sig_logic_x_3 : CKBD0BWP7T port map(I => FE_PHN293_sig_logic_x_3, Z => FE_PHN518_sig_logic_x_3);
  FE_PHC517_sig_logic_y_1 : CKBD0BWP7T port map(I => FE_PHN529_sig_logic_y_1, Z => FE_PHN517_sig_logic_y_1);
  FE_PHC516_sig_logic_y_3 : CKBD0BWP7T port map(I => FE_PHN523_sig_logic_y_3, Z => FE_PHN516_sig_logic_y_3);
  FE_PHC515_gl_ram_n_1111 : DEL01BWP7T port map(I => FE_PHN515_gl_ram_n_1111, Z => FE_PHN277_gl_ram_n_1111);
  FE_PHC514_sig_logic_x_2 : CKBD2BWP7T port map(I => FE_PHN514_sig_logic_x_2, Z => FE_PHN455_sig_logic_x_2);
  FE_PHC513_sig_logic_x_0 : CKBD0BWP7T port map(I => FE_PHN513_sig_logic_x_0, Z => sig_logic_x(0));
  FE_PHC512_sig_logic_x_1 : BUFFD0BWP7T port map(I => FE_PHN512_sig_logic_x_1, Z => FE_PHN506_sig_logic_x_1);
  FE_PHC511_ml_ms_tb_n_5 : DEL01BWP7T port map(I => ml_ms_tb_n_5, Z => FE_PHN511_ml_ms_tb_n_5);
  FE_PHC510_gl_ram_n_1111 : CKBD0BWP7T port map(I => FE_PHN510_gl_ram_n_1111, Z => FE_PHN487_gl_ram_n_1111);
  FE_PHC509_ml_ms_tb_n_5 : CKBD0BWP7T port map(I => FE_PHN511_ml_ms_tb_n_5, Z => FE_PHN509_ml_ms_tb_n_5);
  FE_PHC508_ml_ms_cnt_n_7 : DEL01BWP7T port map(I => ml_ms_cnt_n_7, Z => FE_PHN508_ml_ms_cnt_n_7);
  FE_PHC507_ml_ms_cnt_n_9 : BUFFD3BWP7T port map(I => ml_ms_cnt_n_9, Z => FE_PHN507_ml_ms_cnt_n_9);
  FE_PHC506_sig_logic_x_1 : DEL02BWP7T port map(I => FE_PHN506_sig_logic_x_1, Z => sig_logic_x(1));
  FE_PHC505_sig_logic_x_0 : DEL02BWP7T port map(I => sig_logic_x(0), Z => FE_PHN505_sig_logic_x_0);
  FE_PHC504_ml_ms_count15k_1 : DEL01BWP7T port map(I => FE_PHN504_ml_ms_count15k_1, Z => FE_PHN428_ml_ms_count15k_1);
  FE_PHC503_ml_ms_count25M_3 : DEL0BWP7T port map(I => FE_PHN503_ml_ms_count25M_3, Z => FE_PHN434_ml_ms_count25M_3);
  FE_PHC502_ml_ms_cnt_count_1 : DEL0BWP7T port map(I => ml_ms_cnt_count(1), Z => FE_PHN502_ml_ms_cnt_count_1);
  FE_PHC501_clk15k_in : DEL0BWP7T port map(I => clk15k_in, Z => FE_PHN501_clk15k_in);
  FE_PHC500_ml_ms_cntD_n_22 : DEL1BWP7T port map(I => ml_ms_cntD_n_22, Z => FE_PHN500_ml_ms_cntD_n_22);
  FE_PHC499_ml_ms_cntD_n_12 : DEL1BWP7T port map(I => FE_PHN499_ml_ms_cntD_n_12, Z => ml_ms_cntD_n_12);
  FE_PHC498_ml_ms_cntD_n_13 : DEL1BWP7T port map(I => ml_ms_cntD_n_13, Z => FE_PHN498_ml_ms_cntD_n_13);
  FE_PHC497_ml_il_x1_input_register_3 : DEL1BWP7T port map(I => ml_il_x1_input_register(3), Z => FE_PHN497_ml_il_x1_input_register_3);
  FE_PHC496_ml_ms_cnt_n_17 : DEL1BWP7T port map(I => ml_ms_cnt_n_17, Z => FE_PHN496_ml_ms_cnt_n_17);
  FE_PHC495_ml_ms_cnt_n_15 : DEL1BWP7T port map(I => ml_ms_cnt_n_15, Z => FE_PHN495_ml_ms_cnt_n_15);
  FE_PHC494_ml_ms_cnt_n_21 : DEL1BWP7T port map(I => FE_PHN494_ml_ms_cnt_n_21, Z => ml_ms_cnt_n_21);
  FE_PHC493_ml_ms_cnt_n_22 : DEL1BWP7T port map(I => ml_ms_cnt_n_22, Z => FE_PHN493_ml_ms_cnt_n_22);
  FE_PHC492_ml_ms_cnt_n_19 : DEL1BWP7T port map(I => ml_ms_cnt_n_19, Z => FE_PHN492_ml_ms_cnt_n_19);
  FE_PHC491_ml_ms_cntD_n_9 : DEL1BWP7T port map(I => ml_ms_cntD_n_9, Z => FE_PHN491_ml_ms_cntD_n_9);
  FE_PHC490_ml_ms_cntD_n_11 : DEL1BWP7T port map(I => FE_PHN490_ml_ms_cntD_n_11, Z => ml_ms_cntD_n_11);
  FE_PHC489_ml_ms_cntD_n_10 : DEL1BWP7T port map(I => ml_ms_cntD_n_10, Z => FE_PHN489_ml_ms_cntD_n_10);
  FE_PHC488_ml_ms_ed_n_8 : DEL1BWP7T port map(I => ml_ms_ed_n_8, Z => FE_PHN488_ml_ms_ed_n_8);
  FE_PHC487_gl_ram_n_1111 : DEL0BWP7T port map(I => FE_PHN487_gl_ram_n_1111, Z => FE_PHN283_gl_ram_n_1111);
  FE_PHC486_ml_ms_btnflipfloprst : DEL1BWP7T port map(I => FE_PHN486_ml_ms_btnflipfloprst, Z => ml_ms_btnflipfloprst);
  FE_PHC485_ml_il_y1_n_47 : DEL0BWP7T port map(I => ml_il_y1_n_47, Z => FE_PHN485_ml_il_y1_n_47);
  FE_PHC484_ml_il_x1_n_47 : DEL0BWP7T port map(I => ml_il_x1_n_47, Z => FE_PHN484_ml_il_x1_n_47);
  FE_PHC483_ml_il_y1_input_register_3 : DEL1BWP7T port map(I => ml_il_y1_input_register(3), Z => FE_PHN483_ml_il_y1_input_register_3);
  FE_PHC482_ml_il_y1_n_48 : DEL0BWP7T port map(I => ml_il_y1_n_48, Z => FE_PHN482_ml_il_y1_n_48);
  FE_PHC481_ml_il_x1_n_48 : DEL0BWP7T port map(I => ml_il_x1_n_48, Z => FE_PHN481_ml_il_x1_n_48);
  FE_PHC480_ml_ms_n_58 : DEL1BWP7T port map(I => ml_ms_n_58, Z => FE_PHN480_ml_ms_n_58);
  FE_PHC479_ml_il_y1_n_49 : CKBD0BWP7T port map(I => ml_il_y1_n_49, Z => FE_PHN479_ml_il_y1_n_49);
  FE_PHC478_ml_ms_mfsm_n_46 : DEL1BWP7T port map(I => FE_PHN478_ml_ms_mfsm_n_46, Z => ml_ms_mfsm_n_46);
  FE_PHC477_ml_ms_mfsm_n_45 : DEL1BWP7T port map(I => ml_ms_mfsm_n_45, Z => FE_PHN477_ml_ms_mfsm_n_45);
  FE_PHC476_ml_ms_mfsm_n_43 : DEL1BWP7T port map(I => ml_ms_mfsm_n_43, Z => FE_PHN476_ml_ms_mfsm_n_43);
  FE_PHC475_ml_ms_tb_n_6 : DEL1BWP7T port map(I => FE_PHN475_ml_ms_tb_n_6, Z => ml_ms_tb_n_6);
  FE_PHC474_ml_ms_cnt_n_11 : DEL1BWP7T port map(I => FE_PHN474_ml_ms_cnt_n_11, Z => ml_ms_cnt_n_11);
  FE_PHC473_ml_ms_mfsm_n_29 : DEL1BWP7T port map(I => FE_PHN473_ml_ms_mfsm_n_29, Z => ml_ms_mfsm_n_29);
  FE_PHC472_ml_ms_cnt_n_10 : DEL0BWP7T port map(I => ml_ms_cnt_n_10, Z => FE_PHN472_ml_ms_cnt_n_10);
  FE_PHC471_ml_ms_n_57 : DEL1BWP7T port map(I => ml_ms_n_57, Z => FE_PHN471_ml_ms_n_57);
  FE_PHC470_ml_ms_n_54 : DEL1BWP7T port map(I => ml_ms_n_54, Z => FE_PHN470_ml_ms_n_54);
  FE_PHC469_ml_ms_n_60 : DEL1BWP7T port map(I => ml_ms_n_60, Z => FE_PHN469_ml_ms_n_60);
  FE_PHC468_gl_vgd_n_64 : DEL1BWP7T port map(I => gl_vgd_n_64, Z => FE_PHN468_gl_vgd_n_64);
  FE_PHC467_ml_ms_ed_n_2 : DEL1BWP7T port map(I => ml_ms_ed_n_2, Z => FE_PHN467_ml_ms_ed_n_2);
  FE_PHC466_ml_ms_mfsm_n_42 : DEL1BWP7T port map(I => FE_PHN466_ml_ms_mfsm_n_42, Z => ml_ms_mfsm_n_42);
  FE_PHC465_ml_ms_n_25 : DEL1BWP7T port map(I => FE_PHN465_ml_ms_n_25, Z => ml_ms_n_25);
  FE_PHC464_ml_ms_n_34 : DEL1BWP7T port map(I => FE_PHN464_ml_ms_n_34, Z => ml_ms_n_34);
  FE_PHC463_ml_ms_n_31 : DEL1BWP7T port map(I => ml_ms_n_31, Z => FE_PHN463_ml_ms_n_31);
  FE_PHC462_ml_ms_n_24 : DEL1BWP7T port map(I => ml_ms_n_24, Z => FE_PHN462_ml_ms_n_24);
  FE_PHC461_ml_ms_n_26 : DEL1BWP7T port map(I => FE_PHN461_ml_ms_n_26, Z => ml_ms_n_26);
  FE_PHC460_ml_ms_n_30 : DEL1BWP7T port map(I => ml_ms_n_30, Z => FE_PHN460_ml_ms_n_30);
  FE_PHC459_ml_ms_n_20 : DEL1BWP7T port map(I => FE_PHN459_ml_ms_n_20, Z => ml_ms_n_20);
  FE_PHC458_ml_ms_n_32 : DEL1BWP7T port map(I => ml_ms_n_32, Z => FE_PHN458_ml_ms_n_32);
  FE_PHC457_ml_ms_n_19 : DEL1BWP7T port map(I => FE_PHN457_ml_ms_n_19, Z => ml_ms_n_19);
  FE_PHC456_ml_ms_ed_n_5 : DEL1BWP7T port map(I => FE_PHN456_ml_ms_ed_n_5, Z => ml_ms_ed_n_5);
  FE_PHC455_sig_logic_x_2 : DEL0BWP7T port map(I => FE_PHN455_sig_logic_x_2, Z => sig_logic_x(2));
  FE_PHC454_ml_ms_mfsm_state_0 : DEL1BWP7T port map(I => ml_ms_mfsm_state(0), Z => FE_PHN454_ml_ms_mfsm_state_0);
  FE_PHC453_gl_vgd_horizontal_counter_7 : DEL1BWP7T port map(I => FE_PHN453_gl_vgd_horizontal_counter_7, Z => gl_vgd_horizontal_counter(7));
  FE_PHC452_ml_ms_mfsm_n_47 : DEL0BWP7T port map(I => FE_PHN452_ml_ms_mfsm_n_47, Z => ml_ms_mfsm_n_47);
  FE_PHC451_gl_vgd_horizontal_counter_8 : DEL1BWP7T port map(I => gl_vgd_horizontal_counter(8), Z => FE_PHN451_gl_vgd_horizontal_counter_8);
  FE_PHC450_gl_vgd_horizontal_counter_6 : DEL1BWP7T port map(I => gl_vgd_horizontal_counter(6), Z => FE_PHN450_gl_vgd_horizontal_counter_6);
  FE_PHC449_gl_vgd_horizontal_counter_4 : DEL1BWP7T port map(I => gl_vgd_horizontal_counter(4), Z => FE_PHN449_gl_vgd_horizontal_counter_4);
  FE_PHC448_gl_vgd_horizontal_counter_2 : DEL2BWP7T port map(I => gl_vgd_horizontal_counter(2), Z => FE_PHN448_gl_vgd_horizontal_counter_2);
  FE_PHC447_ml_ms_cnt_count_1 : DEL02BWP7T port map(I => FE_PHN502_ml_ms_cnt_count_1, Z => FE_PHN447_ml_ms_cnt_count_1);
  FE_PHC446_gl_vgd_horizontal_counter_5 : DEL3BWP7T port map(I => gl_vgd_horizontal_counter(5), Z => FE_PHN446_gl_vgd_horizontal_counter_5);
  FE_PHC445_gl_vgd_horizontal_counter_3 : DEL1BWP7T port map(I => gl_vgd_horizontal_counter(3), Z => FE_PHN445_gl_vgd_horizontal_counter_3);
  FE_PHC444_gl_vgd_horizontal_counter_1 : DEL1BWP7T port map(I => FE_PHN444_gl_vgd_horizontal_counter_1, Z => gl_vgd_horizontal_counter(1));
  FE_PHC443_ml_ms_mfsm_state_2 : DEL02BWP7T port map(I => FE_PHN443_ml_ms_mfsm_state_2, Z => ml_ms_mfsm_state(2));
  FE_PHC442_gl_vgd_vertical_counter_9 : DEL1BWP7T port map(I => FE_PHN442_gl_vgd_vertical_counter_9, Z => gl_vgd_vertical_counter(9));
  FE_PHC441_ml_il_x1_state_0 : DEL1BWP7T port map(I => ml_il_x1_state(0), Z => FE_PHN441_ml_il_x1_state_0);
  FE_PHC440_ml_buttons_mouse_0 : DEL1BWP7T port map(I => FE_PHN440_ml_buttons_mouse_0, Z => ml_buttons_mouse(0));
  FE_PHC439_ml_ms_count25M_5 : DEL02BWP7T port map(I => FE_PHN439_ml_ms_count25M_5, Z => ml_ms_count25M(5));
  FE_PHC438_clk15k_in : DEL02BWP7T port map(I => FE_PHN501_clk15k_in, Z => FE_PHN438_clk15k_in);
  FE_PHC437_ml_ms_count25M_4 : DEL0BWP7T port map(I => ml_ms_count25M(4), Z => FE_PHN437_ml_ms_count25M_4);
  FE_PHC436_ml_ms_count25M_7 : DEL1BWP7T port map(I => FE_PHN436_ml_ms_count25M_7, Z => ml_ms_count25M(7));
  FE_PHC435_gl_vgd_horizontal_counter_0 : DEL1BWP7T port map(I => FE_PHN435_gl_vgd_horizontal_counter_0, Z => gl_vgd_horizontal_counter(0));
  FE_PHC434_ml_ms_count25M_3 : DEL02BWP7T port map(I => FE_PHN434_ml_ms_count25M_3, Z => ml_ms_count25M(3));
  FE_PHC433_gl_vgd_vertical_counter_7 : DEL1BWP7T port map(I => FE_PHN433_gl_vgd_vertical_counter_7, Z => gl_vgd_vertical_counter(7));
  FE_PHC432_gl_vgd_horizontal_counter_9 : DEL1BWP7T port map(I => FE_PHN432_gl_vgd_horizontal_counter_9, Z => gl_vgd_horizontal_counter(9));
  FE_PHC431_ml_il_x1_state_1 : DEL1BWP7T port map(I => FE_PHN431_ml_il_x1_state_1, Z => ml_il_x1_state(1));
  FE_PHC430_gl_gr_lg_lv_n_11 : DEL1BWP7T port map(I => gl_gr_lg_lv_n_11, Z => FE_PHN430_gl_gr_lg_lv_n_11);
  FE_PHC429_ml_mouseX_2 : DEL1BWP7T port map(I => FE_PHN429_ml_mouseX_2, Z => ml_mouseX(2));
  FE_PHC428_ml_ms_count15k_1 : DEL0BWP7T port map(I => FE_PHN428_ml_ms_count15k_1, Z => ml_ms_count15k(1));
  FE_PHC427_ml_ms_count25M_10 : DEL1BWP7T port map(I => FE_PHN427_ml_ms_count25M_10, Z => ml_ms_count25M(10));
  FE_PHC426_gl_gr_lg_lv_n_10 : DEL0BWP7T port map(I => gl_gr_lg_lv_n_10, Z => FE_PHN426_gl_gr_lg_lv_n_10);
  FE_PHC425_ml_ms_mux_select : DEL1BWP7T port map(I => ml_ms_mux_select, Z => FE_PHN425_ml_ms_mux_select);
  FE_PHC424_ml_il_y1_state_0 : DEL1BWP7T port map(I => ml_il_y1_state(0), Z => FE_PHN424_ml_il_y1_state_0);
  FE_PHC423_gl_vgd_vertical_counter_5 : DEL1BWP7T port map(I => FE_PHN423_gl_vgd_vertical_counter_5, Z => gl_vgd_vertical_counter(5));
  FE_PHC422_ml_ms_count15k_2 : DEL02BWP7T port map(I => ml_ms_count15k(2), Z => FE_PHN422_ml_ms_count15k_2);
  FE_PHC421_gl_vgd_vertical_counter_6 : DEL1BWP7T port map(I => FE_PHN421_gl_vgd_vertical_counter_6, Z => gl_vgd_vertical_counter(6));
  FE_PHC420_ml_buttons_mouse_1 : DEL1BWP7T port map(I => ml_buttons_mouse(1), Z => FE_PHN420_ml_buttons_mouse_1);
  FE_PHC419_gl_vgd_vertical_counter_3 : DEL2BWP7T port map(I => gl_vgd_vertical_counter(3), Z => FE_PHN419_gl_vgd_vertical_counter_3);
  FE_PHC418_gl_vgd_vertical_counter_4 : DEL1BWP7T port map(I => FE_PHN418_gl_vgd_vertical_counter_4, Z => gl_vgd_vertical_counter(4));
  FE_PHC417_ml_ms_count15k_3 : DEL0BWP7T port map(I => ml_ms_count15k(3), Z => FE_PHN417_ml_ms_count15k_3);
  FE_PHC416_ml_ms_sfsm_state_0 : DEL1BWP7T port map(I => ml_ms_sfsm_state(0), Z => FE_PHN416_ml_ms_sfsm_state_0);
  FE_PHC415_ml_ms_count25M_6 : DEL1BWP7T port map(I => ml_ms_count25M(6), Z => FE_PHN415_ml_ms_count25M_6);
  FE_PHC414_ml_ms_count15k_0 : DEL1BWP7T port map(I => FE_PHN414_ml_ms_count15k_0, Z => ml_ms_count15k(0));
  FE_PHC413_gl_sig_scale_h : DEL2BWP7T port map(I => gl_sig_scale_h, Z => FE_PHN413_gl_sig_scale_h);
  FE_PHC412_gl_vgd_vertical_counter_0 : DEL1BWP7T port map(I => gl_vgd_vertical_counter(0), Z => FE_PHN412_gl_vgd_vertical_counter_0);
  FE_PHC411_ml_ms_data_sr_11bit_7 : DEL1BWP7T port map(I => ml_ms_data_sr_11bit(7), Z => FE_PHN411_ml_ms_data_sr_11bit_7);
  FE_PHC410_gl_vgd_vertical_counter_1 : DEL1BWP7T port map(I => FE_PHN410_gl_vgd_vertical_counter_1, Z => gl_vgd_vertical_counter(1));
  FE_PHC409_gl_vgd_vertical_counter_2 : DEL1BWP7T port map(I => gl_vgd_vertical_counter(2), Z => FE_PHN409_gl_vgd_vertical_counter_2);
  FE_PHC408_ml_ms_count25M_2 : DEL1BWP7T port map(I => FE_PHN408_ml_ms_count25M_2, Z => ml_ms_count25M(2));
  FE_PHC407_gl_gr_lg_lh_n_9 : DEL1BWP7T port map(I => gl_gr_lg_lh_n_9, Z => FE_PHN407_gl_gr_lg_lh_n_9);
  FE_PHC406_gl_gr_lg_lh_n_14 : DEL1BWP7T port map(I => gl_gr_lg_lh_n_14, Z => FE_PHN406_gl_gr_lg_lh_n_14);
  FE_PHC405_gl_gr_lg_lv_n_14 : DEL1BWP7T port map(I => gl_gr_lg_lv_n_14, Z => FE_PHN405_gl_gr_lg_lv_n_14);
  FE_PHC404_data_in : DEL1BWP7T port map(I => data_in, Z => FE_PHN404_data_in);
  FE_PHC403_gl_gr_lg_lh_n_11 : DEL1BWP7T port map(I => FE_PHN403_gl_gr_lg_lh_n_11, Z => gl_gr_lg_lh_n_11);
  FE_PHC402_ml_il_y1_state_1 : DEL1BWP7T port map(I => ml_il_y1_state(1), Z => FE_PHN402_ml_il_y1_state_1);
  FE_PHC401_ml_mouseY_0 : DEL1BWP7T port map(I => ml_mouseY(0), Z => FE_PHN401_ml_mouseY_0);
  FE_PHC400_gl_gr_lg_lv_n_13 : DEL1BWP7T port map(I => FE_PHN400_gl_gr_lg_lv_n_13, Z => gl_gr_lg_lv_n_13);
  FE_PHC399_ml_ms_cntD_count_1 : DEL1BWP7T port map(I => ml_ms_cntD_count(1), Z => FE_PHN399_ml_ms_cntD_count_1);
  FE_PHC398_ml_mouseX_0 : DEL1BWP7T port map(I => ml_mouseX(0), Z => FE_PHN398_ml_mouseX_0);
  FE_PHC397_ml_ms_cntD_n_0 : DEL1BWP7T port map(I => ml_ms_cntD_n_0, Z => FE_PHN397_ml_ms_cntD_n_0);
  FE_PHC396_ml_ms_cnt_n_0 : DEL1BWP7T port map(I => ml_ms_cnt_n_0, Z => FE_PHN396_ml_ms_cnt_n_0);
  FE_PHC395_ml_mouseY_1 : DEL1BWP7T port map(I => ml_mouseY(1), Z => FE_PHN395_ml_mouseY_1);
  FE_PHC394_ml_buttons_mouse_2 : DEL1BWP7T port map(I => ml_buttons_mouse(2), Z => FE_PHN394_ml_buttons_mouse_2);
  FE_PHC393_ml_ms_cntD_n_23 : DEL1BWP7T port map(I => ml_ms_cntD_n_23, Z => FE_PHN393_ml_ms_cntD_n_23);
  FE_PHC392_ml_mouseY_2 : DEL1BWP7T port map(I => ml_mouseY(2), Z => FE_PHN392_ml_mouseY_2);
  FE_PHC391_ml_mouseX_1 : DEL1BWP7T port map(I => ml_mouseX(1), Z => FE_PHN391_ml_mouseX_1);
  FE_PHC390_ml_ms_sr11_data_out_1_80 : DEL1BWP7T port map(I => ml_ms_sr11_data_out_1_80, Z => FE_PHN390_ml_ms_sr11_data_out_1_80);
  FE_PHC389_gl_gr_lg_lh_n_15 : DEL1BWP7T port map(I => gl_gr_lg_lh_n_15, Z => FE_PHN389_gl_gr_lg_lh_n_15);
  FE_PHC388_ml_ms_sr11_data_out_5_84 : DEL1BWP7T port map(I => FE_PHN388_ml_ms_sr11_data_out_5_84, Z => ml_ms_sr11_data_out_5_84);
  FE_PHC387_ml_ms_sr11_data_out_0_79 : DEL1BWP7T port map(I => ml_ms_sr11_data_out_0_79, Z => FE_PHN387_ml_ms_sr11_data_out_0_79);
  FE_PHC386_ml_ms_data_sr_11bit_2 : DEL1BWP7T port map(I => FE_PHN386_ml_ms_data_sr_11bit_2, Z => ml_ms_data_sr_11bit(2));
  FE_PHC385_ml_ms_data_sr_11bit_4 : DEL1BWP7T port map(I => FE_PHN385_ml_ms_data_sr_11bit_4, Z => ml_ms_data_sr_11bit(4));
  FE_PHC384_ml_ms_count_debounce_11 : DEL1BWP7T port map(I => FE_PHN384_ml_ms_count_debounce_11, Z => ml_ms_count_debounce(11));
  FE_PHC383_ml_ms_data_sr_11bit_6 : DEL1BWP7T port map(I => FE_PHN383_ml_ms_data_sr_11bit_6, Z => ml_ms_data_sr_11bit(6));
  FE_PHC382_gl_sig_scale_v : DEL1BWP7T port map(I => gl_sig_scale_v, Z => FE_PHN382_gl_sig_scale_v);
  FE_PHC381_ml_buttons_mouse_4 : DEL2BWP7T port map(I => ml_buttons_mouse(4), Z => FE_PHN381_ml_buttons_mouse_4);
  FE_PHC380_ml_ms_data_sr_11bit_3 : DEL1BWP7T port map(I => FE_PHN380_ml_ms_data_sr_11bit_3, Z => ml_ms_data_sr_11bit(3));
  FE_PHC379_ml_ms_count_debounce_10 : DEL1BWP7T port map(I => FE_PHN379_ml_ms_count_debounce_10, Z => ml_ms_count_debounce(10));
  FE_PHC378_ml_ms_cnt_count_0 : DEL1BWP7T port map(I => FE_PHN378_ml_ms_cnt_count_0, Z => ml_ms_cnt_count(0));
  FE_PHC377_ml_ms_count_debounce_3 : DEL1BWP7T port map(I => ml_ms_count_debounce(3), Z => FE_PHN377_ml_ms_count_debounce_3);
  FE_PHC376_gl_gr_lg_le_new_count_e_1 : DEL2BWP7T port map(I => FE_PHN376_gl_gr_lg_le_new_count_e_1, Z => gl_gr_lg_le_new_count_e(1));
  FE_PHC375_ml_ms_count_debounce_4 : DEL1BWP7T port map(I => ml_ms_count_debounce(4), Z => FE_PHN375_ml_ms_count_debounce_4);
  FE_PHC374_gl_gr_lg_le_new_count_e_6 : DEL2BWP7T port map(I => gl_gr_lg_le_new_count_e(6), Z => FE_PHN374_gl_gr_lg_le_new_count_e_6);
  FE_PHC373_gl_gr_lg_le_new_count_e_8 : DEL2BWP7T port map(I => gl_gr_lg_le_new_count_e(8), Z => FE_PHN373_gl_gr_lg_le_new_count_e_8);
  FE_PHC372_gl_gr_lg_le_new_count_e_9 : DEL2BWP7T port map(I => gl_gr_lg_le_new_count_e(9), Z => FE_PHN372_gl_gr_lg_le_new_count_e_9);
  FE_PHC371_gl_gr_lg_le_new_count_e_7 : DEL2BWP7T port map(I => gl_gr_lg_le_new_count_e(7), Z => FE_PHN371_gl_gr_lg_le_new_count_e_7);
  FE_PHC370_ml_ms_ed_reg1 : DEL1BWP7T port map(I => FE_PHN370_ml_ms_ed_reg1, Z => ml_ms_ed_reg1);
  FE_PHC369_gl_gr_lg_le_new_count_e_5 : DEL2BWP7T port map(I => gl_gr_lg_le_new_count_e(5), Z => FE_PHN369_gl_gr_lg_le_new_count_e_5);
  FE_PHC368_gl_gr_lg_lv_l_edge_reg1 : DEL1BWP7T port map(I => gl_gr_lg_lv_l_edge_reg1, Z => FE_PHN368_gl_gr_lg_lv_l_edge_reg1);
  FE_PHC367_gl_gr_lg_le_new_count_e_0 : DEL2BWP7T port map(I => gl_gr_lg_le_new_count_e(0), Z => FE_PHN367_gl_gr_lg_le_new_count_e_0);
  FE_PHC366_gl_gr_lg_le_new_count_e_3 : DEL2BWP7T port map(I => gl_gr_lg_le_new_count_e(3), Z => FE_PHN366_gl_gr_lg_le_new_count_e_3);
  FE_PHC365_gl_gr_lg_lh_l_edge_reg1 : DEL1BWP7T port map(I => gl_gr_lg_lh_l_edge_reg1, Z => FE_PHN365_gl_gr_lg_lh_l_edge_reg1);
  FE_PHC364_gl_gr_lg_le_new_count_e_4 : DEL2BWP7T port map(I => gl_gr_lg_le_new_count_e(4), Z => FE_PHN364_gl_gr_lg_le_new_count_e_4);
  FE_PHC363_gl_gr_lg_le_new_count_e_2 : DEL2BWP7T port map(I => gl_gr_lg_le_new_count_e(2), Z => FE_PHN363_gl_gr_lg_le_new_count_e_2);
  FE_PHC362_ml_ms_ed_state_1 : DEL1BWP7T port map(I => FE_PHN362_ml_ms_ed_state_1, Z => ml_ms_ed_state(1));
  FE_PHC361_ml_ms_count_debounce_9 : DEL1BWP7T port map(I => ml_ms_count_debounce(9), Z => FE_PHN361_ml_ms_count_debounce_9);
  FE_PHC360_ml_ms_count_debounce_8 : DEL1BWP7T port map(I => ml_ms_count_debounce(8), Z => FE_PHN360_ml_ms_count_debounce_8);
  FE_PHC359_gl_vgd_vertical_counter_8 : DEL1BWP7T port map(I => FE_PHN359_gl_vgd_vertical_counter_8, Z => gl_vgd_vertical_counter(8));
  FE_PHC358_ml_buttons_mouse_3 : DEL1BWP7T port map(I => ml_buttons_mouse(3), Z => FE_PHN358_ml_buttons_mouse_3);
  FE_PHC357_ml_ms_cntD_count_0 : DEL1BWP7T port map(I => FE_PHN357_ml_ms_cntD_count_0, Z => ml_ms_cntD_count(0));
  FE_PHC356_ml_ms_cntD_count_2 : DEL1BWP7T port map(I => ml_ms_cntD_count(2), Z => FE_PHN356_ml_ms_cntD_count_2);
  FE_PSC355_gl_ram_ram_16_2 : BUFFD1BWP7T port map(I => gl_ram_ram_16(2), Z => FE_PSN355_gl_ram_ram_16_2);
  FE_PSC354_gl_ram_ram_73_2 : BUFFD1BWP7T port map(I => gl_ram_ram_73(2), Z => FE_PSN354_gl_ram_ram_73_2);
  FE_PSC353_gl_ram_ram_36_2 : BUFFD1BWP7T port map(I => gl_ram_ram_36(2), Z => FE_PSN353_gl_ram_ram_36_2);
  FE_PSC352_gl_ram_ram_85_2 : BUFFD1BWP7T port map(I => gl_ram_ram_85(2), Z => FE_PSN352_gl_ram_ram_85_2);
  FE_PSC351_gl_ram_ram_72_2 : BUFFD1BWP7T port map(I => gl_ram_ram_72(2), Z => FE_PSN351_gl_ram_ram_72_2);
  FE_PSC350_gl_ram_ram_55_2 : BUFFD1BWP7T port map(I => gl_ram_ram_55(2), Z => FE_PSN350_gl_ram_ram_55_2);
  FE_PHC349_FE_OFN4_gl_ram_n_1111 : CKBD0BWP7T port map(I => FE_PHN334_FE_OFN4_gl_ram_n_1111, Z => FE_PHN349_FE_OFN4_gl_ram_n_1111);
  FE_PHC348_FE_OFN4_gl_ram_n_1111 : CKBD0BWP7T port map(I => FE_PHN332_FE_OFN4_gl_ram_n_1111, Z => FE_PHN348_FE_OFN4_gl_ram_n_1111);
  FE_PHC347_FE_OFN4_gl_ram_n_1111 : CKBD0BWP7T port map(I => FE_PHN330_FE_OFN4_gl_ram_n_1111, Z => FE_PHN347_FE_OFN4_gl_ram_n_1111);
  FE_PHC346_FE_OFN4_gl_ram_n_1111 : CKBD1BWP7T port map(I => FE_PHN329_FE_OFN4_gl_ram_n_1111, Z => FE_PHN346_FE_OFN4_gl_ram_n_1111);
  FE_PHC345_FE_OFN4_gl_ram_n_1111 : CKBD1BWP7T port map(I => FE_PHN333_FE_OFN4_gl_ram_n_1111, Z => FE_PHN345_FE_OFN4_gl_ram_n_1111);
  FE_PHC344_FE_OFN4_gl_ram_n_1111 : BUFFD0BWP7T port map(I => FE_PHN326_FE_OFN4_gl_ram_n_1111, Z => FE_PHN344_FE_OFN4_gl_ram_n_1111);
  FE_PHC343_FE_OFN4_gl_ram_n_1111 : CKBD0BWP7T port map(I => FE_PHN328_FE_OFN4_gl_ram_n_1111, Z => FE_PHN343_FE_OFN4_gl_ram_n_1111);
  FE_PHC342_FE_OFN4_gl_ram_n_1111 : CKBD0BWP7T port map(I => FE_PHN327_FE_OFN4_gl_ram_n_1111, Z => FE_PHN342_FE_OFN4_gl_ram_n_1111);
  FE_PHC341_FE_OFN4_gl_ram_n_1111 : DEL01BWP7T port map(I => FE_PHN322_FE_OFN4_gl_ram_n_1111, Z => FE_PHN341_FE_OFN4_gl_ram_n_1111);
  FE_PHC340_FE_OFN4_gl_ram_n_1111 : CKBD0BWP7T port map(I => FE_PHN331_FE_OFN4_gl_ram_n_1111, Z => FE_PHN340_FE_OFN4_gl_ram_n_1111);
  FE_PHC339_FE_OFN4_gl_ram_n_1111 : DEL015BWP7T port map(I => FE_PHN324_FE_OFN4_gl_ram_n_1111, Z => FE_PHN339_FE_OFN4_gl_ram_n_1111);
  FE_PHC338_FE_OFN4_gl_ram_n_1111 : BUFFD0BWP7T port map(I => FE_PHN320_FE_OFN4_gl_ram_n_1111, Z => FE_PHN338_FE_OFN4_gl_ram_n_1111);
  FE_PHC337_FE_OFN4_gl_ram_n_1111 : CKBD0BWP7T port map(I => FE_PHN323_FE_OFN4_gl_ram_n_1111, Z => FE_PHN337_FE_OFN4_gl_ram_n_1111);
  FE_PHC336_FE_OFN4_gl_ram_n_1111 : DEL01BWP7T port map(I => FE_PHN321_FE_OFN4_gl_ram_n_1111, Z => FE_PHN336_FE_OFN4_gl_ram_n_1111);
  FE_PHC335_FE_OFN4_gl_ram_n_1111 : BUFFD1BWP7T port map(I => FE_OFN4_gl_ram_n_1111, Z => FE_PHN335_FE_OFN4_gl_ram_n_1111);
  FE_PHC334_FE_OFN4_gl_ram_n_1111 : BUFFD1BWP7T port map(I => FE_OFN4_gl_ram_n_1111, Z => FE_PHN334_FE_OFN4_gl_ram_n_1111);
  FE_PHC333_FE_OFN4_gl_ram_n_1111 : BUFFD0BWP7T port map(I => FE_OFN4_gl_ram_n_1111, Z => FE_PHN333_FE_OFN4_gl_ram_n_1111);
  FE_PHC332_FE_OFN4_gl_ram_n_1111 : BUFFD1BWP7T port map(I => FE_OFN4_gl_ram_n_1111, Z => FE_PHN332_FE_OFN4_gl_ram_n_1111);
  FE_PHC331_FE_OFN4_gl_ram_n_1111 : CKBD1BWP7T port map(I => FE_OFN4_gl_ram_n_1111, Z => FE_PHN331_FE_OFN4_gl_ram_n_1111);
  FE_PHC330_FE_OFN4_gl_ram_n_1111 : BUFFD1BWP7T port map(I => FE_OFN4_gl_ram_n_1111, Z => FE_PHN330_FE_OFN4_gl_ram_n_1111);
  FE_PHC329_FE_OFN4_gl_ram_n_1111 : BUFFD0BWP7T port map(I => FE_OFN4_gl_ram_n_1111, Z => FE_PHN329_FE_OFN4_gl_ram_n_1111);
  FE_PHC328_FE_OFN4_gl_ram_n_1111 : DEL01BWP7T port map(I => FE_OFN4_gl_ram_n_1111, Z => FE_PHN328_FE_OFN4_gl_ram_n_1111);
  FE_PHC327_FE_OFN4_gl_ram_n_1111 : CKBD2BWP7T port map(I => FE_OFN4_gl_ram_n_1111, Z => FE_PHN327_FE_OFN4_gl_ram_n_1111);
  FE_PHC326_FE_OFN4_gl_ram_n_1111 : CKBD10BWP7T port map(I => FE_OFN4_gl_ram_n_1111, Z => FE_PHN326_FE_OFN4_gl_ram_n_1111);
  FE_PHC325_FE_OFN4_gl_ram_n_1111 : CKBD6BWP7T port map(I => FE_PHN522_FE_OFN4_gl_ram_n_1111, Z => FE_PHN325_FE_OFN4_gl_ram_n_1111);
  FE_PHC324_FE_OFN4_gl_ram_n_1111 : CKBD12BWP7T port map(I => FE_OFN4_gl_ram_n_1111, Z => FE_PHN324_FE_OFN4_gl_ram_n_1111);
  FE_PHC323_FE_OFN4_gl_ram_n_1111 : CKBD12BWP7T port map(I => FE_OFN4_gl_ram_n_1111, Z => FE_PHN323_FE_OFN4_gl_ram_n_1111);
  FE_PHC322_FE_OFN4_gl_ram_n_1111 : CKBD10BWP7T port map(I => FE_OFN4_gl_ram_n_1111, Z => FE_PHN322_FE_OFN4_gl_ram_n_1111);
  FE_PHC321_FE_OFN4_gl_ram_n_1111 : CKBD12BWP7T port map(I => FE_OFN4_gl_ram_n_1111, Z => FE_PHN321_FE_OFN4_gl_ram_n_1111);
  FE_PHC320_FE_OFN4_gl_ram_n_1111 : CKBD12BWP7T port map(I => FE_OFN4_gl_ram_n_1111, Z => FE_PHN320_FE_OFN4_gl_ram_n_1111);
  FE_PHC319_gl_ram_n_1111 : BUFFD0BWP7T port map(I => FE_PHN308_gl_ram_n_1111, Z => FE_PHN319_gl_ram_n_1111);
  FE_PHC318_gl_ram_n_1111 : BUFFD0BWP7T port map(I => FE_PHN313_gl_ram_n_1111, Z => FE_PHN318_gl_ram_n_1111);
  FE_PHC317_gl_ram_n_1111 : CKBD1BWP7T port map(I => FE_PHN301_gl_ram_n_1111, Z => FE_PHN317_gl_ram_n_1111);
  FE_PHC316_sig_logic_y_3 : BUFFD4BWP7T port map(I => sig_logic_y(3), Z => FE_PHN316_sig_logic_y_3);
  FE_PHC315_sig_logic_x_2 : DEL01BWP7T port map(I => sig_logic_x(2), Z => FE_PHN315_sig_logic_x_2);
  FE_PHC314_sig_logic_x_3 : CKBD0BWP7T port map(I => FE_PHN518_sig_logic_x_3, Z => FE_PHN314_sig_logic_x_3);
  FE_PHC313_gl_ram_n_1111 : BUFFD0BWP7T port map(I => FE_PHN307_gl_ram_n_1111, Z => FE_PHN313_gl_ram_n_1111);
  FE_PHC312_gl_ram_n_1111 : BUFFD0BWP7T port map(I => FE_PHN298_gl_ram_n_1111, Z => FE_PHN312_gl_ram_n_1111);
  FE_PHC311_gl_ram_n_1111 : BUFFD0BWP7T port map(I => FE_PHN312_gl_ram_n_1111, Z => FE_PHN311_gl_ram_n_1111);
  FE_PHC310_gl_ram_n_1111 : DEL0BWP7T port map(I => FE_PHN298_gl_ram_n_1111, Z => FE_PHN310_gl_ram_n_1111);
  FE_PHC309_gl_ram_n_1111 : DEL0BWP7T port map(I => FE_PHN318_gl_ram_n_1111, Z => FE_PHN309_gl_ram_n_1111);
  FE_PHC308_gl_ram_n_1111 : BUFFD1BWP7T port map(I => FE_PHN311_gl_ram_n_1111, Z => FE_PHN308_gl_ram_n_1111);
  FE_PHC307_gl_ram_n_1111 : BUFFD0BWP7T port map(I => FE_PHN520_gl_ram_n_1111, Z => FE_PHN307_gl_ram_n_1111);
  FE_PHC306_gl_ram_n_1111 : BUFFD0BWP7T port map(I => FE_PHN298_gl_ram_n_1111, Z => FE_PHN306_gl_ram_n_1111);
  FE_PHC305_gl_ram_n_1111 : DEL0BWP7T port map(I => FE_PHN319_gl_ram_n_1111, Z => FE_PHN305_gl_ram_n_1111);
  FE_PHC304_gl_ram_n_1111 : BUFFD0BWP7T port map(I => FE_PHN306_gl_ram_n_1111, Z => FE_PHN304_gl_ram_n_1111);
  FE_PHC303_gl_ram_n_1111 : DEL1BWP7T port map(I => FE_PHN298_gl_ram_n_1111, Z => FE_PHN303_gl_ram_n_1111);
  FE_PHC302_gl_ram_n_1111 : BUFFD4BWP7T port map(I => FE_PHN298_gl_ram_n_1111, Z => FE_PHN302_gl_ram_n_1111);
  FE_PHC301_gl_ram_n_1111 : DEL0BWP7T port map(I => FE_PHN310_gl_ram_n_1111, Z => FE_PHN521_gl_ram_n_1111);
  FE_PHC300_gl_ram_n_1111 : DEL1BWP7T port map(I => FE_PHN302_gl_ram_n_1111, Z => FE_PHN300_gl_ram_n_1111);
  FE_PHC299_gl_ram_n_1111 : CKBD2BWP7T port map(I => FE_PHN301_gl_ram_n_1111, Z => FE_PHN299_gl_ram_n_1111);
  FE_PHC298_gl_ram_n_1111 : CKBD12BWP7T port map(I => FE_PHN297_gl_ram_n_1111, Z => FE_PHN298_gl_ram_n_1111);
  FE_PHC297_gl_ram_n_1111 : CKBD12BWP7T port map(I => FE_PHN288_gl_ram_n_1111, Z => FE_PHN297_gl_ram_n_1111);
  FE_PHC296_gl_ram_n_1310 : CKBD0BWP7T port map(I => FE_PHN284_gl_ram_n_1310, Z => FE_PHN296_gl_ram_n_1310);
  FE_PHC295_gl_ram_n_1111 : CKBD0BWP7T port map(I => FE_PHN283_gl_ram_n_1111, Z => FE_PHN295_gl_ram_n_1111);
  FE_PHC294_gl_ram_n_1311 : CKBD0BWP7T port map(I => gl_ram_n_1311, Z => FE_PHN294_gl_ram_n_1311);
  FE_PHC293_sig_logic_x_3 : CKBD0BWP7T port map(I => FE_PHN527_sig_logic_x_3, Z => FE_PHN293_sig_logic_x_3);
  FE_PHC292_gl_ram_n_819 : DEL0BWP7T port map(I => FE_PHN519_gl_ram_n_819, Z => FE_PHN292_gl_ram_n_819);
  FE_PHC291_gl_ram_n_1310 : DEL02BWP7T port map(I => FE_PHN296_gl_ram_n_1310, Z => FE_PHN291_gl_ram_n_1310);
  FE_PHC290_gl_ram_n_1111 : CKBD0BWP7T port map(I => FE_PHN295_gl_ram_n_1111, Z => FE_PHN290_gl_ram_n_1111);
  FE_PHC289_gl_ram_n_1111 : DEL02BWP7T port map(I => FE_PHN304_gl_ram_n_1111, Z => FE_PHN289_gl_ram_n_1111);
  FE_PHC288_gl_ram_n_1111 : DEL015BWP7T port map(I => FE_PHN276_gl_ram_n_1111, Z => FE_PHN288_gl_ram_n_1111);
  FE_PHC287_sig_logic_x_3 : CKBD0BWP7T port map(I => sig_logic_x(3), Z => FE_PHN287_sig_logic_x_3);
  FE_PHC286_sig_logic_x_2 : DEL0BWP7T port map(I => FE_PHN315_sig_logic_x_2, Z => FE_PHN286_sig_logic_x_2);
  FE_PHC285_gl_ram_n_819 : DEL0BWP7T port map(I => gl_ram_n_819, Z => FE_PHN285_gl_ram_n_819);
  FE_PHC284_gl_ram_n_1310 : DEL0BWP7T port map(I => gl_ram_n_1310, Z => FE_PHN284_gl_ram_n_1310);
  FE_PHC283_gl_ram_n_1111 : DEL0BWP7T port map(I => FE_PHN280_gl_ram_n_1111, Z => FE_PHN510_gl_ram_n_1111);
  FE_PHC282_gl_ram_n_1111 : DEL1BWP7T port map(I => FE_PHN277_gl_ram_n_1111, Z => FE_PHN282_gl_ram_n_1111);
  FE_PHC281_gl_ram_n_1111 : DEL4BWP7T port map(I => FE_PHN282_gl_ram_n_1111, Z => FE_PHN281_gl_ram_n_1111);
  FE_PHC280_gl_ram_n_1111 : DEL4BWP7T port map(I => FE_PHN278_gl_ram_n_1111, Z => FE_PHN280_gl_ram_n_1111);
  FE_PHC279_gl_ram_n_1111 : DEL4BWP7T port map(I => FE_PHN281_gl_ram_n_1111, Z => FE_PHN279_gl_ram_n_1111);
  FE_PHC278_gl_ram_n_1111 : DEL4BWP7T port map(I => FE_PHN279_gl_ram_n_1111, Z => FE_PHN278_gl_ram_n_1111);
  FE_PHC277_gl_ram_n_1111 : DEL4BWP7T port map(I => gl_ram_n_1111, Z => FE_PHN515_gl_ram_n_1111);
  FE_PHC276_gl_ram_n_1111 : DEL4BWP7T port map(I => FE_PHN290_gl_ram_n_1111, Z => FE_PHN276_gl_ram_n_1111);
  FE_OCPC275_gl_ram_ram_9_0 : BUFFD1BWP7T port map(I => gl_ram_ram_9(0), Z => FE_OCPN275_gl_ram_ram_9_0);
  FE_OCPC274_gl_ram_ram_32_1 : BUFFD1BWP7T port map(I => gl_ram_ram_32(1), Z => FE_OCPN274_gl_ram_ram_32_1);
  FE_OCPC273_gl_ram_ram_13_2 : BUFFD1BWP7T port map(I => gl_ram_ram_13(2), Z => FE_OCPN273_gl_ram_ram_13_2);
  FE_OCPC272_gl_ram_ram_43_0 : BUFFD1BWP7T port map(I => gl_ram_ram_43(0), Z => FE_OCPN272_gl_ram_ram_43_0);
  FE_OCPC271_gl_ram_ram_40_2 : BUFFD1BWP7T port map(I => gl_ram_ram_40(2), Z => FE_OCPN271_gl_ram_ram_40_2);
  FE_OCPC270_gl_ram_ram_24_2 : BUFFD1BWP7T port map(I => gl_ram_ram_24(2), Z => FE_OCPN270_gl_ram_ram_24_2);
  FE_OCPC269_gl_ram_ram_52_0 : BUFFD1BWP7T port map(I => gl_ram_ram_52(0), Z => FE_OCPN269_gl_ram_ram_52_0);
  FE_RC_207_0 : INVD1BWP7T port map(I => gl_ram_n_90, ZN => FE_RN_89_0);
  FE_RC_206_0 : IND2D2BWP7T port map(A1 => FE_RN_89_0, B1 => gl_ram_ram_69(0), ZN => FE_RN_90_0);
  FE_RC_205_0 : ND2D2BWP7T port map(A1 => gl_ram_n_265, A2 => FE_RN_90_0, ZN => gl_ram_n_1498);
  FE_OCPC268_gl_ram_ram_10_0 : BUFFD1BWP7T port map(I => gl_ram_ram_10(0), Z => FE_OCPN268_gl_ram_ram_10_0);
  FE_OCPC267_gl_ram_ram_63_0 : BUFFD1BWP7T port map(I => gl_ram_ram_63(0), Z => FE_OCPN267_gl_ram_ram_63_0);
  FE_OCPC266_gl_ram_ram_55_0 : BUFFD1BWP7T port map(I => gl_ram_ram_55(0), Z => FE_OCPN266_gl_ram_ram_55_0);
  FE_RC_204_0 : ND2D3BWP7T port map(A1 => gl_ram_ram_56(1), A2 => gl_ram_n_89, ZN => FE_RN_88_0);
  FE_RC_203_0 : IOA21D2BWP7T port map(A1 => gl_ram_ram_59(1), A2 => gl_ram_n_87, B => FE_RN_88_0, ZN => gl_ram_n_1539);
  FE_RC_202_0 : ND2D2BWP7T port map(A1 => gl_ram_ram_88(0), A2 => gl_ram_n_89, ZN => FE_RN_87_0);
  FE_RC_201_0 : ND2D2BWP7T port map(A1 => gl_ram_n_235, A2 => FE_RN_87_0, ZN => gl_ram_n_1504);
  FE_RC_200_0 : ND2D2BWP7T port map(A1 => gl_ram_ram_6(2), A2 => gl_ram_n_93, ZN => FE_RN_86_0);
  FE_RC_199_0 : ND2D2BWP7T port map(A1 => gl_ram_n_274, A2 => FE_RN_86_0, ZN => gl_ram_n_1495);
  FE_RC_198_0 : IND2D2BWP7T port map(A1 => FE_RN_72_0, B1 => gl_ram_ram_49(0), ZN => FE_RN_73_0);
  FE_RC_197_0 : INVD1BWP7T port map(I => gl_ram_n_92, ZN => FE_RN_85_0);
  FE_RC_196_0 : IND2D2BWP7T port map(A1 => FE_RN_85_0, B1 => gl_ram_ram_55(0), ZN => gl_ram_n_209);
  FE_RC_195_0 : IND2D2BWP7T port map(A1 => FE_RN_41_0, B1 => gl_ram_ram_50(0), ZN => gl_ram_n_216);
  FE_OCPC265_gl_ram_ram_54_0 : BUFFD1BWP7T port map(I => gl_ram_ram_54(0), Z => FE_OCPN265_gl_ram_ram_54_0);
  FE_OCPC264_gl_ram_ram_30_0 : BUFFD1BWP7T port map(I => gl_ram_ram_30(0), Z => FE_OCPN264_gl_ram_ram_30_0);
  FE_OCPC263_gl_ram_ram_4_0 : BUFFD1BWP7T port map(I => gl_ram_ram_4(0), Z => FE_OCPN263_gl_ram_ram_4_0);
  FE_OCPC262_gl_ram_ram_49_0 : BUFFD1BWP7T port map(I => gl_ram_ram_49(0), Z => FE_OCPN262_gl_ram_ram_49_0);
  FE_OCPC260_gl_ram_ram_2_0 : BUFFD0BWP7T port map(I => gl_ram_ram_2(0), Z => FE_OCPN260_gl_ram_ram_2_0);
  FE_OCPC259_gl_ram_ram_9_0 : BUFFD0BWP7T port map(I => FE_OCPN275_gl_ram_ram_9_0, Z => FE_OCPN259_gl_ram_ram_9_0);
  FE_OCPC257_gl_ram_ram_42_0 : BUFFD1BWP7T port map(I => gl_ram_ram_42(0), Z => FE_OCPN257_gl_ram_ram_42_0);
  FE_OCPC255_gl_ram_ram_15_0 : BUFFD0BWP7T port map(I => gl_ram_ram_15(0), Z => FE_OCPN255_gl_ram_ram_15_0);
  FE_RC_194_0 : INVD1BWP7T port map(I => gl_ram_n_87, ZN => FE_RN_84_0);
  FE_RC_193_0 : IND2D2BWP7T port map(A1 => FE_RN_84_0, B1 => gl_ram_ram_51(0), ZN => gl_ram_n_176);
  FE_RC_192_0 : ND2D2BWP7T port map(A1 => gl_ram_ram_94(0), A2 => gl_ram_n_93, ZN => FE_RN_83_0);
  FE_RC_191_0 : ND2D2BWP7T port map(A1 => gl_ram_n_239, A2 => FE_RN_83_0, ZN => gl_ram_n_1438);
  FE_RC_190_0 : INVD1BWP7T port map(I => gl_ram_n_89, ZN => FE_RN_81_0);
  FE_RC_189_0 : IND2D2BWP7T port map(A1 => FE_RN_81_0, B1 => gl_ram_ram_40(0), ZN => FE_RN_82_0);
  FE_RC_188_0 : ND2D2BWP7T port map(A1 => gl_ram_n_213, A2 => FE_RN_82_0, ZN => gl_ram_n_1510);
  FE_RC_187_0 : INVD1BWP7T port map(I => gl_ram_n_86, ZN => FE_RN_80_0);
  FE_RC_186_0 : IND2D2BWP7T port map(A1 => FE_RN_80_0, B1 => gl_ram_ram_42(0), ZN => gl_ram_n_215);
  FE_RC_185_0 : IND2D2BWP7T port map(A1 => FE_RN_39_0, B1 => gl_ram_ram_54(0), ZN => FE_RN_40_0);
  FE_RC_184_0 : IND2D2BWP7T port map(A1 => FE_RN_37_0, B1 => gl_ram_ram_52(0), ZN => FE_RN_38_0);
  FE_RC_183_0 : AOI21D2BWP7T port map(A1 => gl_ram_n_582, A2 => gl_ram_n_581, B => gl_ram_n_97, ZN => gl_ram_n_684);
  FE_RC_182_0 : CKND2BWP7T port map(I => gl_ram_n_89, ZN => FE_RN_78_0);
  FE_RC_181_0 : IND2D2BWP7T port map(A1 => FE_RN_78_0, B1 => gl_ram_ram_32(2), ZN => FE_RN_79_0);
  FE_RC_180_0 : ND2D2BWP7T port map(A1 => gl_ram_n_305, A2 => FE_RN_79_0, ZN => gl_ram_n_1487);
  FE_OCPC252_gl_ram_ram_25_2 : BUFFD1BWP7T port map(I => gl_ram_ram_25(2), Z => FE_OCPN252_gl_ram_ram_25_2);
  FE_OCPC250_gl_ram_ram_24_2 : BUFFD1BWP7T port map(I => FE_OCPN270_gl_ram_ram_24_2, Z => FE_OCPN250_gl_ram_ram_24_2);
  FE_OCPC249_gl_ram_ram_48_2 : BUFFD1BWP7T port map(I => gl_ram_ram_48(2), Z => FE_OCPN249_gl_ram_ram_48_2);
  FE_OCPC248_gl_ram_ram_51_2 : BUFFD1BWP7T port map(I => gl_ram_ram_51(2), Z => FE_OCPN248_gl_ram_ram_51_2);
  FE_OCPC247_gl_ram_ram_41_2 : BUFFD1BWP7T port map(I => gl_ram_ram_41(2), Z => FE_OCPN247_gl_ram_ram_41_2);
  FE_OCPC246_gl_ram_ram_1_2 : BUFFD0BWP7T port map(I => gl_ram_ram_1(2), Z => FE_OCPN246_gl_ram_ram_1_2);
  FE_OCPC245_gl_ram_ram_5_0 : BUFFD1BWP7T port map(I => gl_ram_ram_5(0), Z => FE_OCPN245_gl_ram_ram_5_0);
  FE_OCPC244_gl_ram_ram_29_2 : BUFFD1BWP7T port map(I => gl_ram_ram_29(2), Z => FE_OCPN244_gl_ram_ram_29_2);
  FE_OCPC243_gl_ram_ram_28_0 : BUFFD1BWP7T port map(I => gl_ram_ram_28(0), Z => FE_OCPN243_gl_ram_ram_28_0);
  FE_OCPC242_gl_ram_ram_55_1 : BUFFD1BWP7T port map(I => gl_ram_ram_55(1), Z => FE_OCPN242_gl_ram_ram_55_1);
  FE_RC_179_0 : ND2D1BWP7T port map(A1 => gl_ram_ram_94(2), A2 => gl_ram_n_93, ZN => FE_RN_77_0);
  FE_RC_178_0 : ND2D1BWP7T port map(A1 => gl_ram_n_340, A2 => FE_RN_77_0, ZN => gl_ram_n_1474);
  FE_RC_177_0 : ND2D3BWP7T port map(A1 => gl_ram_n_643, A2 => gl_ram_n_642, ZN => FE_RN_76_0);
  FE_RC_176_0 : CKND2D4BWP7T port map(A1 => FE_RN_76_0, A2 => gl_ram_n_563, ZN => gl_ram_n_671);
  FE_RC_175_0 : CKND2D2BWP7T port map(A1 => gl_ram_ram_37(0), A2 => gl_ram_n_90, ZN => FE_RN_75_0);
  FE_RC_174_0 : IOA21D2BWP7T port map(A1 => gl_ram_ram_39(0), A2 => gl_ram_n_92, B => FE_RN_75_0, ZN => gl_ram_n_1513);
  FE_RC_173_0 : CKND2D2BWP7T port map(A1 => gl_ram_ram_32(0), A2 => gl_ram_n_89, ZN => FE_RN_74_0);
  FE_RC_172_0 : ND2D2BWP7T port map(A1 => FE_RN_74_0, A2 => gl_ram_n_191, ZN => gl_ram_n_1515);
  FE_RC_171_0 : INVD1BWP7T port map(I => gl_ram_n_88, ZN => FE_RN_72_0);
  FE_RC_169_0 : ND2D3BWP7T port map(A1 => FE_RN_73_0, A2 => gl_ram_n_216, ZN => gl_ram_n_1523);
  FE_RC_168_0 : AOI21D2BWP7T port map(A1 => gl_ram_n_1445, A2 => gl_ram_n_599, B => gl_ram_n_99, ZN => gl_ram_n_685);
  FE_RC_167_0 : INVD8BWP7T port map(I => FE_RN_71_0, ZN => gl_ram_n_1449);
  FE_RC_166_0 : AN2D4BWP7T port map(A1 => gl_ram_n_733, A2 => gl_ram_n_728, Z => FE_RN_71_0);
  FE_RC_165_0 : CKND2D2BWP7T port map(A1 => gl_ram_ram_34(0), A2 => gl_ram_n_86, ZN => FE_RN_70_0);
  FE_RC_164_0 : ND2D2P5BWP7T port map(A1 => FE_RN_70_0, A2 => gl_ram_n_194, ZN => gl_ram_n_1516);
  FE_RC_163_0 : ND2D2BWP7T port map(A1 => gl_ram_ram_29(2), A2 => gl_ram_n_90, ZN => FE_RN_69_0);
  FE_RC_162_0 : IOA21D2BWP7T port map(A1 => gl_ram_ram_31(2), A2 => gl_ram_n_92, B => FE_RN_69_0, ZN => gl_ram_n_1483);
  FE_OCPC240_gl_ram_ram_53_2 : BUFFD1BWP7T port map(I => gl_ram_ram_53(2), Z => FE_OCPN240_gl_ram_ram_53_2);
  FE_OCPC239_gl_ram_ram_86_2 : BUFFD1BWP7T port map(I => gl_ram_ram_86(2), Z => FE_OCPN239_gl_ram_ram_86_2);
  FE_OCPC238_gl_ram_ram_69_2 : BUFFD0BWP7T port map(I => gl_ram_ram_69(2), Z => FE_OCPN238_gl_ram_ram_69_2);
  FE_OCPC237_gl_ram_ram_75_2 : BUFFD0BWP7T port map(I => gl_ram_ram_75(2), Z => FE_OCPN237_gl_ram_ram_75_2);
  FE_OCPC236_gl_ram_ram_82_2 : BUFFD1BWP7T port map(I => gl_ram_ram_82(2), Z => FE_OCPN236_gl_ram_ram_82_2);
  FE_OCPC235_gl_ram_ram_73_2 : BUFFD1BWP7T port map(I => FE_PSN354_gl_ram_ram_73_2, Z => FE_OCPN235_gl_ram_ram_73_2);
  FE_OCPC233_gl_ram_ram_12_1 : BUFFD1BWP7T port map(I => gl_ram_ram_12(1), Z => FE_OCPN233_gl_ram_ram_12_1);
  FE_OCPC231_gl_ram_ram_50_2 : BUFFD1BWP7T port map(I => gl_ram_ram_50(2), Z => FE_OCPN231_gl_ram_ram_50_2);
  FE_OCPC228_gl_ram_ram_72_2 : BUFFD1BWP7T port map(I => FE_PSN351_gl_ram_ram_72_2, Z => FE_OCPN228_gl_ram_ram_72_2);
  FE_OCPC226_gl_ram_ram_46_2 : BUFFD1BWP7T port map(I => gl_ram_ram_46(2), Z => FE_OCPN226_gl_ram_ram_46_2);
  FE_OCPC225_gl_ram_ram_80_2 : BUFFD0BWP7T port map(I => gl_ram_ram_80(2), Z => FE_OCPN225_gl_ram_ram_80_2);
  FE_OCPC221_gl_ram_ram_0_2 : BUFFD0BWP7T port map(I => gl_ram_ram_0(2), Z => FE_OCPN221_gl_ram_ram_0_2);
  FE_OCPC219_gl_ram_ram_87_2 : BUFFD1BWP7T port map(I => gl_ram_ram_87(2), Z => FE_OCPN219_gl_ram_ram_87_2);
  FE_OCPC218_gl_ram_ram_71_2 : BUFFD1BWP7T port map(I => gl_ram_ram_71(2), Z => FE_OCPN218_gl_ram_ram_71_2);
  FE_OCPC217_gl_ram_ram_67_2 : BUFFD0BWP7T port map(I => gl_ram_ram_67(2), Z => FE_OCPN217_gl_ram_ram_67_2);
  FE_OCPC214_gl_ram_ram_18_2 : BUFFD0BWP7T port map(I => gl_ram_ram_18(2), Z => FE_OCPN214_gl_ram_ram_18_2);
  FE_OCPC210_gl_ram_ram_12_2 : BUFFD1BWP7T port map(I => gl_ram_ram_12(2), Z => FE_OCPN210_gl_ram_ram_12_2);
  FE_OCPC208_gl_ram_ram_15_2 : BUFFD1BWP7T port map(I => gl_ram_ram_15(2), Z => FE_OCPN208_gl_ram_ram_15_2);
  FE_OCPC204_gl_ram_ram_79_2 : BUFFD1BWP7T port map(I => gl_ram_ram_79(2), Z => FE_OCPN204_gl_ram_ram_79_2);
  FE_OCPC203_gl_ram_ram_44_2 : BUFFD1BWP7T port map(I => gl_ram_ram_44(2), Z => FE_OCPN203_gl_ram_ram_44_2);
  FE_OCPC200_gl_ram_ram_47_2 : BUFFD0BWP7T port map(I => gl_ram_ram_47(2), Z => FE_OCPN200_gl_ram_ram_47_2);
  FE_OCPC199_gl_ram_ram_2_2 : BUFFD1BWP7T port map(I => gl_ram_ram_2(2), Z => FE_OCPN199_gl_ram_ram_2_2);
  FE_OCPC198_gl_ram_ram_65_2 : BUFFD0BWP7T port map(I => gl_ram_ram_65(2), Z => FE_OCPN198_gl_ram_ram_65_2);
  FE_OCPC197_gl_ram_ram_8_2 : BUFFD0BWP7T port map(I => gl_ram_ram_8(2), Z => FE_OCPN197_gl_ram_ram_8_2);
  FE_OCPC196_gl_ram_ram_78_2 : BUFFD1BWP7T port map(I => gl_ram_ram_78(2), Z => FE_OCPN196_gl_ram_ram_78_2);
  FE_OCPC195_gl_ram_ram_23_2 : BUFFD0BWP7T port map(I => gl_ram_ram_23(2), Z => FE_OCPN195_gl_ram_ram_23_2);
  FE_OCPC194_gl_ram_ram_3_2 : BUFFD1BWP7T port map(I => gl_ram_ram_3(2), Z => FE_OCPN194_gl_ram_ram_3_2);
  FE_OCPC193_gl_ram_ram_92_2 : BUFFD1BWP7T port map(I => gl_ram_ram_92(2), Z => FE_OCPN193_gl_ram_ram_92_2);
  FE_OCPC192_gl_ram_ram_77_2 : BUFFD1BWP7T port map(I => gl_ram_ram_77(2), Z => FE_OCPN192_gl_ram_ram_77_2);
  FE_OCPC191_gl_ram_ram_83_2 : BUFFD1BWP7T port map(I => gl_ram_ram_83(2), Z => FE_OCPN191_gl_ram_ram_83_2);
  FE_OCPC189_gl_ram_ram_52_0 : BUFFD0BWP7T port map(I => FE_OCPN269_gl_ram_ram_52_0, Z => FE_OCPN189_gl_ram_ram_52_0);
  FE_OCPC186_gl_ram_ram_13_0 : BUFFD1BWP7T port map(I => gl_ram_ram_13(0), Z => FE_OCPN186_gl_ram_ram_13_0);
  FE_OCPC184_gl_ram_ram_54_1 : BUFFD1BWP7T port map(I => gl_ram_ram_54(1), Z => FE_OCPN184_gl_ram_ram_54_1);
  FE_RC_161_0 : INVD1BWP7T port map(I => gl_ram_n_90, ZN => FE_RN_67_0);
  FE_RC_160_0 : IND2D2BWP7T port map(A1 => FE_RN_67_0, B1 => gl_ram_ram_85(2), ZN => FE_RN_68_0);
  FE_RC_159_0 : ND2D3BWP7T port map(A1 => FE_RN_68_0, A2 => gl_ram_n_351, ZN => gl_ram_n_1470);
  FE_RC_158_0 : CKND2D2BWP7T port map(A1 => gl_ram_ram_73(2), A2 => gl_ram_n_88, ZN => FE_RN_66_0);
  FE_RC_157_0 : IOA21D2BWP7T port map(A1 => gl_ram_ram_74(2), A2 => gl_ram_n_86, B => FE_RN_66_0, ZN => gl_ram_n_1464);
  FE_RC_156_0 : ND2D2BWP7T port map(A1 => gl_ram_ram_86(2), A2 => gl_ram_n_93, ZN => FE_RN_65_0);
  FE_RC_155_0 : ND2D2BWP7T port map(A1 => FE_RN_65_0, A2 => gl_ram_n_346, ZN => gl_ram_n_1471);
  FE_RC_154_0 : INVD1BWP7T port map(I => gl_ram_n_86, ZN => FE_RN_64_0);
  FE_RC_153_0 : IND2D2BWP7T port map(A1 => FE_RN_64_0, B1 => gl_ram_ram_50(1), ZN => gl_ram_n_379);
  FE_RC_152_0 : CKND2D2BWP7T port map(A1 => gl_ram_ram_61(1), A2 => gl_ram_n_90, ZN => FE_RN_63_0);
  FE_RC_151_0 : ND2D3BWP7T port map(A1 => gl_ram_n_146, A2 => FE_RN_63_0, ZN => gl_ram_n_1538);
  FE_RC_150_0 : IOA21D2BWP7T port map(A1 => gl_ram_ram_1(0), A2 => gl_ram_n_88, B => gl_ram_n_173, ZN => gl_ram_n_1525);
  FE_RC_149_0 : ND2D2BWP7T port map(A1 => gl_ram_ram_45(2), A2 => gl_ram_n_90, ZN => FE_RN_62_0);
  FE_RC_148_0 : ND2D3BWP7T port map(A1 => gl_ram_n_326, A2 => FE_RN_62_0, ZN => gl_ram_n_1479);
  FE_OCPC183_gl_ram_ram_5_2 : BUFFD1BWP7T port map(I => gl_ram_ram_5(2), Z => FE_OCPN183_gl_ram_ram_5_2);
  FE_OCPC180_gl_ram_ram_6_2 : BUFFD1BWP7T port map(I => gl_ram_ram_6(2), Z => FE_OCPN180_gl_ram_ram_6_2);
  FE_OCPC179_gl_ram_ram_99_2 : BUFFD1BWP7T port map(I => gl_ram_ram_99(2), Z => FE_OCPN179_gl_ram_ram_99_2);
  FE_RC_147_0 : INVD1BWP7T port map(I => gl_ram_n_90, ZN => FE_RN_60_0);
  FE_RC_146_0 : IND2D2BWP7T port map(A1 => FE_RN_60_0, B1 => gl_ram_ram_61(2), ZN => FE_RN_61_0);
  FE_RC_145_0 : ND2D3BWP7T port map(A1 => gl_ram_n_335, A2 => FE_RN_61_0, ZN => gl_ram_n_1477);
  FE_RC_144_0 : CKND2D2BWP7T port map(A1 => gl_ram_ram_78(2), A2 => gl_ram_n_93, ZN => FE_RN_59_0);
  FE_RC_143_0 : ND2D2BWP7T port map(A1 => FE_RN_59_0, A2 => gl_ram_n_362, ZN => gl_ram_n_1465);
  FE_OCPC175_gl_ram_ram_37_0 : BUFFD1BWP7T port map(I => gl_ram_ram_37(0), Z => FE_OCPN175_gl_ram_ram_37_0);
  FE_RC_142_0 : CKND2D2BWP7T port map(A1 => gl_ram_ram_30(0), A2 => gl_ram_n_93, ZN => FE_RN_58_0);
  FE_RC_141_0 : ND2D2P5BWP7T port map(A1 => FE_RN_58_0, A2 => gl_ram_n_207, ZN => gl_ram_n_459);
  FE_OCPC174_gl_ram_ram_0_1 : BUFFD0BWP7T port map(I => gl_ram_ram_0(1), Z => FE_OCPN174_gl_ram_ram_0_1);
  FE_OCPC173_gl_ram_ram_7_2 : BUFFD0BWP7T port map(I => gl_ram_ram_7(2), Z => FE_OCPN173_gl_ram_ram_7_2);
  FE_RC_140_0 : CKND2D3BWP7T port map(A1 => gl_ram_ram_30(2), A2 => gl_ram_n_93, ZN => FE_RN_57_0);
  FE_RC_139_0 : ND2D3BWP7T port map(A1 => FE_RN_57_0, A2 => gl_ram_n_316, ZN => gl_ram_n_510);
  FE_RC_138_0 : AOI21D2BWP7T port map(A1 => gl_ram_n_650, A2 => gl_ram_n_631, B => gl_ram_n_96, ZN => gl_ram_n_683);
  FE_RC_137_0 : INVD1BWP7T port map(I => gl_ram_n_91, ZN => FE_RN_56_0);
  FE_RC_136_0 : IND2D2BWP7T port map(A1 => FE_RN_56_0, B1 => gl_ram_ram_44(2), ZN => gl_ram_n_324);
  FE_RC_135_0 : ND2D3BWP7T port map(A1 => gl_ram_n_614, A2 => gl_ram_n_615, ZN => FE_RN_55_0);
  FE_RC_134_0 : ND2D4BWP7T port map(A1 => FE_RN_55_0, A2 => FE_RN_24_0, ZN => gl_ram_n_8);
  FE_RC_133_0 : INVD2BWP7T port map(I => gl_ram_ram_97(2), ZN => FE_RN_54_0);
  FE_RC_132_0 : NR2XD1BWP7T port map(A1 => FE_RN_54_0, A2 => gl_ram_n_259, ZN => gl_ram_n_3);
  FE_RC_131_0 : INVD1BWP7T port map(I => gl_ram_n_93, ZN => FE_RN_52_0);
  FE_RC_130_0 : IND2D2BWP7T port map(A1 => FE_RN_52_0, B1 => gl_ram_ram_46(2), ZN => FE_RN_53_0);
  FE_RC_129_0 : ND2D3BWP7T port map(A1 => FE_RN_53_0, A2 => gl_ram_n_324, ZN => gl_ram_n_1480);
  FE_RC_128_0 : ND2D2BWP7T port map(A1 => gl_ram_ram_53(0), A2 => gl_ram_n_90, ZN => FE_RN_51_0);
  FE_RC_127_0 : ND2D2BWP7T port map(A1 => gl_ram_n_209, A2 => FE_RN_51_0, ZN => gl_ram_n_1512);
  FE_RC_126_0 : ND2D2BWP7T port map(A1 => gl_ram_ram_0(0), A2 => gl_ram_n_89, ZN => FE_RN_50_0);
  FE_RC_125_0 : ND2D2BWP7T port map(A1 => gl_ram_n_171, A2 => FE_RN_50_0, ZN => gl_ram_n_1505);
  FE_RC_124_0 : CKND2D2BWP7T port map(A1 => gl_ram_ram_46(1), A2 => gl_ram_n_93, ZN => FE_RN_49_0);
  FE_RC_123_0 : ND2D3BWP7T port map(A1 => FE_RN_49_0, A2 => gl_ram_n_135, ZN => gl_ram_n_1541);
  FE_RC_122_0 : INVD1BWP7T port map(I => gl_ram_n_93, ZN => FE_RN_47_0);
  FE_RC_121_0 : IND2D2BWP7T port map(A1 => FE_RN_47_0, B1 => gl_ram_ram_6(0), ZN => FE_RN_48_0);
  FE_RC_120_0 : ND2D2BWP7T port map(A1 => gl_ram_n_162, A2 => FE_RN_48_0, ZN => gl_ram_n_1506);
  FE_RC_119_0 : INVD1BWP7T port map(I => gl_ram_n_89, ZN => FE_RN_45_0);
  FE_RC_118_0 : IND2D2BWP7T port map(A1 => FE_RN_45_0, B1 => gl_ram_ram_48(0), ZN => FE_RN_46_0);
  FE_RC_117_0 : ND2D2BWP7T port map(A1 => gl_ram_n_176, A2 => FE_RN_46_0, ZN => gl_ram_n_1524);
  FE_RC_116_0 : ND2D2BWP7T port map(A1 => gl_ram_ram_5(1), A2 => gl_ram_n_90, ZN => FE_RN_44_0);
  FE_RC_115_0 : IOA21D2BWP7T port map(A1 => gl_ram_ram_7(1), A2 => gl_ram_n_92, B => FE_RN_44_0, ZN => gl_ram_n_1459);
  FE_RC_114_0 : ND2D2BWP7T port map(A1 => gl_ram_ram_40(2), A2 => gl_ram_n_89, ZN => FE_RN_43_0);
  FE_RC_113_0 : IOA21D2BWP7T port map(A1 => gl_ram_ram_43(2), A2 => gl_ram_n_87, B => FE_RN_43_0, ZN => gl_ram_n_1482);
  FE_RC_112_0 : CKND2D2BWP7T port map(A1 => gl_ram_ram_9(1), A2 => gl_ram_n_88, ZN => FE_RN_42_0);
  FE_RC_111_0 : ND2D2BWP7T port map(A1 => FE_RN_42_0, A2 => gl_ram_n_398, ZN => gl_ram_n_1454);
  FE_OCPC170_gl_ram_ram_40_0 : BUFFD1BWP7T port map(I => gl_ram_ram_40(0), Z => FE_OCPN170_gl_ram_ram_40_0);
  FE_OCPC169_gl_ram_ram_57_2 : BUFFD1BWP7T port map(I => gl_ram_ram_57(2), Z => FE_OCPN169_gl_ram_ram_57_2);
  FE_OCPC167_gl_ram_n_14 : BUFFD1BWP7T port map(I => gl_ram_n_14, Z => FE_OCPN167_gl_ram_n_14);
  FE_RC_110_0 : INVD1BWP7T port map(I => gl_ram_n_86, ZN => FE_RN_41_0);
  FE_RC_108_0 : INVD1BWP7T port map(I => gl_ram_n_91, ZN => FE_RN_37_0);
  FE_RC_106_0 : INVD1BWP7T port map(I => gl_ram_n_93, ZN => FE_RN_39_0);
  FE_RC_104_0 : ND2D3BWP7T port map(A1 => FE_RN_40_0, A2 => FE_RN_38_0, ZN => gl_ram_n_1522);
  FE_RC_102_0 : AOI21D2BWP7T port map(A1 => gl_ram_n_604, A2 => gl_ram_n_602, B => gl_ram_n_94, ZN => gl_ram_n_688);
  FE_RC_99_0 : ND2D2BWP7T port map(A1 => gl_ram_ram_27(2), A2 => gl_ram_n_87, ZN => FE_RN_35_0);
  FE_RC_98_0 : ND2D2BWP7T port map(A1 => FE_RN_35_0, A2 => gl_ram_n_350, ZN => gl_ram_n_508);
  FE_OCPC163_gl_ram_ram_21_2 : BUFFD1BWP7T port map(I => gl_ram_ram_21(2), Z => FE_OCPN163_gl_ram_ram_21_2);
  FE_RC_97_0 : INVD1BWP7T port map(I => gl_ram_n_92, ZN => FE_RN_32_0);
  FE_RC_96_0 : IND2D2BWP7T port map(A1 => FE_RN_32_0, B1 => gl_ram_ram_55(1), ZN => FE_RN_33_0);
  FE_RC_95_0 : IND2D2BWP7T port map(A1 => FE_RN_13_0, B1 => gl_ram_ram_53(1), ZN => FE_RN_34_0);
  FE_RC_94_0 : ND2D2BWP7T port map(A1 => FE_RN_34_0, A2 => FE_RN_33_0, ZN => gl_ram_n_543);
  FE_RC_93_0 : INVD1BWP7T port map(I => gl_ram_n_562, ZN => FE_RN_30_0);
  FE_RC_92_0 : ND2D2BWP7T port map(A1 => gl_ram_n_622, A2 => gl_ram_n_625, ZN => FE_RN_31_0);
  FE_RC_91_0 : CKND2D4BWP7T port map(A1 => FE_RN_31_0, A2 => FE_RN_30_0, ZN => FE_RN_28_0);
  FE_RC_90_0 : ND2D2BWP7T port map(A1 => gl_ram_ram_46(0), A2 => gl_ram_n_93, ZN => FE_RN_29_0);
  FE_RC_89_0 : ND2D2BWP7T port map(A1 => FE_RN_29_0, A2 => gl_ram_n_218, ZN => gl_ram_n_1509);
  FE_RC_88_0 : AOI21D2BWP7T port map(A1 => gl_ram_n_597, A2 => gl_ram_n_596, B => gl_ram_n_4, ZN => gl_ram_n_693);
  FE_RC_85_0 : ND2D6BWP7T port map(A1 => FE_RN_28_0, A2 => gl_ram_n_9, ZN => gl_ram_n_700);
  FE_RC_84_0 : INVD1BWP7T port map(I => gl_ram_n_557, ZN => FE_RN_26_0);
  FE_RC_83_0 : ND2D2BWP7T port map(A1 => gl_ram_n_616, A2 => gl_ram_n_617, ZN => FE_RN_27_0);
  FE_RC_82_0 : ND2D3BWP7T port map(A1 => FE_RN_27_0, A2 => FE_RN_26_0, ZN => gl_ram_n_9);
  FE_RC_81_0 : AOI21D2BWP7T port map(A1 => gl_ram_n_605, A2 => gl_ram_n_603, B => gl_ram_n_97, ZN => gl_ram_n_686);
  FE_RC_80_0 : AOI21D2BWP7T port map(A1 => gl_ram_n_595, A2 => gl_ram_n_594, B => gl_ram_n_98, ZN => gl_ram_n_673);
  FE_OCPC41_gl_ram_ram_98_2 : CKND1BWP7T port map(I => FE_OCPN167_gl_ram_n_14, ZN => FE_OCPN38_gl_ram_ram_98_2);
  FE_OCPC40_gl_ram_ram_98_2 : INVD2BWP7T port map(I => gl_ram_ram_98(2), ZN => gl_ram_n_14);
  FE_RC_79_0 : AOI21D2BWP7T port map(A1 => gl_ram_n_647, A2 => gl_ram_n_646, B => gl_ram_n_4, ZN => gl_ram_n_696);
  FE_RC_78_0 : CKND1BWP7T port map(I => gl_ram_n_556, ZN => FE_RN_24_0);
  FE_OCPC39_gl_ram_ram_97_1 : CKND1BWP7T port map(I => gl_ram_n_15, ZN => FE_OCPN37_gl_ram_ram_97_1);
  FE_OCPC38_gl_ram_ram_97_1 : INVD3BWP7T port map(I => gl_ram_ram_97(1), ZN => gl_ram_n_15);
  FE_RC_75_0 : AOI21D2BWP7T port map(A1 => gl_ram_n_658, A2 => gl_ram_n_573, B => gl_ram_n_256, ZN => gl_ram_n_714);
  FE_OCPC37_gl_ram_ram_98_0 : CKND1BWP7T port map(I => gl_ram_n_20, ZN => FE_OCPN36_gl_ram_ram_98_0);
  FE_OCPC36_gl_ram_ram_98_0 : INVD4BWP7T port map(I => gl_ram_ram_98(0), ZN => gl_ram_n_20);
  FE_OFC35_V : BUFFD5BWP7T port map(I => FE_OFN35_V, Z => V);
  FE_OFC34_H : BUFFD5BWP7T port map(I => FE_OFN34_H, Z => H);
  FE_OFC33_clk15k_switch : BUFFD5BWP7T port map(I => FE_OFN33_clk15k_switch, Z => clk15k_switch);
  FE_OFC32_logic_1_1_net : DEL01BWP7T port map(I => logic_1_1_net, Z => FE_OFN32_logic_1_1_net);
  FE_OFC31_reset : DEL01BWP7T port map(I => reset, Z => FE_OFN31_reset);
  FE_OFC30_gl_rom_n_18 : BUFFD1P5BWP7T port map(I => FE_OFN29_gl_rom_n_18, Z => FE_OFN30_gl_rom_n_18);
  FE_OFC29_gl_rom_n_18 : BUFFD1P5BWP7T port map(I => FE_OFN28_gl_rom_n_18, Z => FE_OFN29_gl_rom_n_18);
  FE_OFC28_gl_rom_n_18 : BUFFD1P5BWP7T port map(I => gl_rom_n_18, Z => FE_OFN28_gl_rom_n_18);
  FE_OFC27_gl_rom_n_21 : BUFFD1P5BWP7T port map(I => FE_OFN26_gl_rom_n_21, Z => FE_OFN27_gl_rom_n_21);
  FE_OFC26_gl_rom_n_21 : BUFFD2BWP7T port map(I => FE_OFN25_gl_rom_n_21, Z => FE_OFN26_gl_rom_n_21);
  FE_OFC25_gl_rom_n_21 : BUFFD1P5BWP7T port map(I => gl_rom_n_21, Z => FE_OFN25_gl_rom_n_21);
  FE_OFC24_gl_rom_n_20 : BUFFD1P5BWP7T port map(I => FE_OFN23_gl_rom_n_20, Z => FE_OFN24_gl_rom_n_20);
  FE_OFC23_gl_rom_n_20 : BUFFD1P5BWP7T port map(I => FE_OFN22_gl_rom_n_20, Z => FE_OFN23_gl_rom_n_20);
  FE_OFC22_gl_rom_n_20 : CKBD1BWP7T port map(I => gl_rom_n_20, Z => FE_OFN22_gl_rom_n_20);
  FE_OFC21_gl_rom_n_16 : BUFFD1P5BWP7T port map(I => FE_OFN20_gl_rom_n_16, Z => FE_OFN21_gl_rom_n_16);
  FE_OFC20_gl_rom_n_16 : CKND2BWP7T port map(I => FE_OFN18_gl_rom_n_16, ZN => FE_OFN20_gl_rom_n_16);
  FE_OFC19_gl_rom_n_16 : INVD1BWP7T port map(I => FE_OFN18_gl_rom_n_16, ZN => FE_OFN19_gl_rom_n_16);
  FE_OFC18_gl_rom_n_16 : INVD1BWP7T port map(I => gl_rom_n_16, ZN => FE_OFN18_gl_rom_n_16);
  FE_OFC17_gl_rom_n_16 : BUFFD1P5BWP7T port map(I => gl_rom_n_16, Z => FE_OFN17_gl_rom_n_16);
  FE_OFC16_gl_rom_n_22 : BUFFD1P5BWP7T port map(I => FE_OFN15_gl_rom_n_22, Z => FE_OFN16_gl_rom_n_22);
  FE_OFC15_gl_rom_n_22 : BUFFD2BWP7T port map(I => gl_rom_n_22, Z => FE_OFN15_gl_rom_n_22);
  FE_OFC14_gl_rom_n_22 : BUFFD1P5BWP7T port map(I => gl_rom_n_22, Z => FE_OFN14_gl_rom_n_22);
  FE_OFC13_gl_rom_n_19 : BUFFD2BWP7T port map(I => FE_OFN12_gl_rom_n_19, Z => FE_OFN13_gl_rom_n_19);
  FE_OFC12_gl_rom_n_19 : BUFFD2BWP7T port map(I => FE_OFN11_gl_rom_n_19, Z => FE_OFN12_gl_rom_n_19);
  FE_OFC11_gl_rom_n_19 : BUFFD2BWP7T port map(I => gl_rom_n_19, Z => FE_OFN11_gl_rom_n_19);
  FE_OFC10_gl_rom_n_17 : BUFFD1P5BWP7T port map(I => FE_OFN8_gl_rom_n_17, Z => FE_OFN10_gl_rom_n_17);
  FE_OFC9_gl_rom_n_17 : BUFFD1P5BWP7T port map(I => FE_OFN8_gl_rom_n_17, Z => FE_OFN9_gl_rom_n_17);
  FE_OFC8_gl_rom_n_17 : BUFFD2BWP7T port map(I => gl_rom_n_17, Z => FE_OFN8_gl_rom_n_17);
  FE_OFC7_gl_rom_n_15 : BUFFD1P5BWP7T port map(I => FE_OFN6_gl_rom_n_15, Z => FE_OFN7_gl_rom_n_15);
  FE_OFC6_gl_rom_n_15 : BUFFD2BWP7T port map(I => FE_OFN5_gl_rom_n_15, Z => FE_OFN6_gl_rom_n_15);
  FE_OFC5_gl_rom_n_15 : BUFFD2BWP7T port map(I => gl_rom_n_15, Z => FE_OFN5_gl_rom_n_15);
  FE_OFC4_gl_ram_n_1111 : BUFFD2BWP7T port map(I => FE_PHN298_gl_ram_n_1111, Z => FE_OFN4_gl_ram_n_1111);
  CTS_ccl_a_BUF_clk_G0_L5_47 : CKBD0BWP7T port map(I => CTS_363, Z => CTS_362);
  CTS_cex_INV_clk_G0_L5_46 : CKND4BWP7T port map(I => CTS_363, ZN => CTS_361);
  CTS_ccl_a_BUF_clk_G0_L4_20 : CKBD2BWP7T port map(I => gl_ram_n_74, Z => CTS_363);
  CTS_ccl_a_BUF_clk_G0_L5_45 : CKBD0BWP7T port map(I => CTS_360, Z => CTS_359);
  CTS_cex_INV_clk_G0_L5_44 : CKND0BWP7T port map(I => CTS_360, ZN => CTS_358);
  CTS_ccl_a_BUF_clk_G0_L4_19 : CKBD0BWP7T port map(I => gl_ram_n_72, Z => CTS_360);
  CTS_ccl_a_BUF_clk_G0_L5_43 : CKBD0BWP7T port map(I => CTS_357, Z => CTS_356);
  CTS_cex_INV_clk_G0_L5_42 : CKND0BWP7T port map(I => CTS_357, ZN => CTS_355);
  CTS_ccl_a_BUF_clk_G0_L4_18 : CKBD2BWP7T port map(I => gl_ram_n_54, Z => CTS_357);
  CTS_ccl_a_BUF_clk_G0_L5_41 : CKBD0BWP7T port map(I => CTS_354, Z => CTS_353);
  CTS_cex_INV_clk_G0_L5_40 : CKND0BWP7T port map(I => CTS_354, ZN => CTS_352);
  CTS_ccl_a_BUF_clk_G0_L4_17 : CKBD0BWP7T port map(I => gl_ram_n_46, Z => CTS_354);
  CTS_ccl_a_BUF_clk_G0_L5_39 : CKBD0BWP7T port map(I => CTS_351, Z => CTS_350);
  CTS_cex_INV_clk_G0_L5_38 : CKND0BWP7T port map(I => CTS_351, ZN => CTS_349);
  CTS_ccl_a_BUF_clk_G0_L4_16 : CKBD0BWP7T port map(I => gl_ram_n_44, Z => CTS_351);
  CTS_ccl_a_BUF_clk_G0_L5_37 : CKBD4BWP7T port map(I => CTS_348, Z => CTS_347);
  CTS_cex_INV_clk_G0_L5_36 : CKND3BWP7T port map(I => CTS_348, ZN => CTS_346);
  CTS_ccl_a_BUF_clk_G0_L4_15 : CKBD1BWP7T port map(I => gl_ram_n_40, Z => CTS_348);
  CTS_cfo_BUF_clk_G0_L2_3 : CKBD12BWP7T port map(I => CTS_365, Z => CTS_364);
  CTS_ccl_a_BUF_clk_G0_L5_35 : CKBD0BWP7T port map(I => gl_ram_n_103, Z => CTS_343);
  CTS_cex_INV_clk_G0_L5_34 : CKND0BWP7T port map(I => gl_ram_n_103, ZN => CTS_342);
  CTS_ccl_a_BUF_clk_G0_L5_33 : CKBD0BWP7T port map(I => gl_ram_n_101, Z => CTS_341);
  CTS_cex_INV_clk_G0_L5_32 : CKND0BWP7T port map(I => gl_ram_n_101, ZN => CTS_340);
  CTS_ccl_a_BUF_clk_G0_L5_31 : CKBD0BWP7T port map(I => gl_ram_n_84, Z => CTS_339);
  CTS_cex_INV_clk_G0_L5_30 : CKND0BWP7T port map(I => gl_ram_n_84, ZN => CTS_338);
  CTS_ccl_a_BUF_clk_G0_L5_29 : CKBD0BWP7T port map(I => gl_ram_n_80, Z => CTS_337);
  CTS_cex_INV_clk_G0_L5_28 : CKND0BWP7T port map(I => gl_ram_n_80, ZN => CTS_336);
  CTS_ccl_a_BUF_clk_G0_L5_27 : CKBD0BWP7T port map(I => gl_ram_n_76, Z => CTS_335);
  CTS_cex_INV_clk_G0_L5_26 : CKND0BWP7T port map(I => gl_ram_n_76, ZN => CTS_334);
  CTS_ccl_a_BUF_clk_G0_L5_25 : CKBD2BWP7T port map(I => gl_ram_n_60, Z => CTS_333);
  CTS_cex_INV_clk_G0_L5_24 : CKND2BWP7T port map(I => gl_ram_n_60, ZN => CTS_332);
  CTS_ccl_a_BUF_clk_G0_L5_23 : CKBD0BWP7T port map(I => gl_ram_n_50, Z => CTS_331);
  CTS_cex_INV_clk_G0_L5_22 : CKND0BWP7T port map(I => gl_ram_n_50, ZN => CTS_330);
  CTS_ccl_a_BUF_clk_G0_L5_21 : CKBD6BWP7T port map(I => gl_ram_n_48, Z => CTS_329);
  CTS_cex_INV_clk_G0_L5_20 : CKND0BWP7T port map(I => gl_ram_n_48, ZN => CTS_328);
  CTS_ccl_a_BUF_clk_G0_L5_19 : CKBD0BWP7T port map(I => gl_ram_n_42, Z => CTS_327);
  CTS_cex_INV_clk_G0_L5_18 : CKND0BWP7T port map(I => gl_ram_n_42, ZN => CTS_326);
  CTS_ccl_a_BUF_clk_G0_L5_17 : CKBD0BWP7T port map(I => gl_ram_n_38, Z => CTS_325);
  CTS_cex_INV_clk_G0_L5_16 : CKND0BWP7T port map(I => gl_ram_n_38, ZN => CTS_324);
  CTS_cfo_BUF_clk_G0_L3_4 : CKBD12BWP7T port map(I => CTS_345, Z => CTS_344);
  CTS_ccl_a_BUF_clk_G0_L4_14 : CKBD6BWP7T port map(I => CTS_323, Z => CTS_322);
  CTS_ccl_a_BUF_clk_G0_L3_3 : CKBD0BWP7T port map(I => CTS_345, Z => CTS_323);
  CTS_ccl_a_BUF_clk_G0_L5_15 : CKBD0BWP7T port map(I => CTS_321, Z => CTS_320);
  CTS_cex_INV_clk_G0_L5_14 : CKND0BWP7T port map(I => CTS_321, ZN => CTS_319);
  CTS_cid_BUF_clk_G0_L4_13 : CKBD2BWP7T port map(I => gl_ram_n_105, Z => CTS_321);
  CTS_ccl_a_BUF_clk_G0_L6_6 : CKBD2BWP7T port map(I => CTS_317, Z => CTS_316);
  CTS_cex_INV_clk_G0_L6_5 : CKND3BWP7T port map(I => CTS_317, ZN => CTS_315);
  CTS_ccl_a_BUF_clk_G0_L5_13 : CKBD4BWP7T port map(I => CTS_318, Z => CTS_317);
  CTS_cid_BUF_clk_G0_L4_12 : CKBD2BWP7T port map(I => gl_ram_n_82, Z => CTS_318);
  CTS_ccl_a_BUF_clk_G0_L5_12 : CKBD0BWP7T port map(I => CTS_314, Z => CTS_313);
  CTS_cex_INV_clk_G0_L5_11 : CKND8BWP7T port map(I => CTS_314, ZN => CTS_312);
  CTS_cid_BUF_clk_G0_L4_11 : CKBD2BWP7T port map(I => gl_ram_n_78, Z => CTS_314);
  CTS_ccl_a_BUF_clk_G0_L5_10 : CKBD0BWP7T port map(I => CTS_311, Z => CTS_310);
  CTS_cex_INV_clk_G0_L5_9 : CKND0BWP7T port map(I => CTS_311, ZN => CTS_309);
  CTS_cid_BUF_clk_G0_L4_10 : CKBD2BWP7T port map(I => gl_ram_n_70, Z => CTS_311);
  CTS_ccl_a_BUF_clk_G0_L5_8 : CKBD0BWP7T port map(I => CTS_308, Z => CTS_307);
  CTS_cex_INV_clk_G0_L5_7 : CKND1BWP7T port map(I => CTS_308, ZN => CTS_306);
  CTS_cid_BUF_clk_G0_L4_9 : CKBD2BWP7T port map(I => gl_ram_n_68, Z => CTS_308);
  CTS_ccl_a_BUF_clk_G0_L6_4 : CKBD2BWP7T port map(I => CTS_304, Z => CTS_303);
  CTS_cex_INV_clk_G0_L6_3 : CKND2BWP7T port map(I => CTS_304, ZN => CTS_302);
  CTS_ccl_a_BUF_clk_G0_L5_6 : CKBD3BWP7T port map(I => CTS_305, Z => CTS_304);
  CTS_cid_BUF_clk_G0_L4_8 : CKBD2BWP7T port map(I => gl_ram_n_66, Z => CTS_305);
  CTS_ccl_a_BUF_clk_G0_L5_5 : CKBD0BWP7T port map(I => CTS_301, Z => CTS_300);
  CTS_cex_INV_clk_G0_L5_4 : CKND1BWP7T port map(I => CTS_301, ZN => CTS_299);
  CTS_cid_BUF_clk_G0_L4_7 : CKBD2BWP7T port map(I => gl_ram_n_64, Z => CTS_301);
  CTS_ccl_a_BUF_clk_G0_L4_6 : CKBD0BWP7T port map(I => gl_ram_n_58, Z => CTS_298);
  CTS_cex_INV_clk_G0_L4_5 : CKND0BWP7T port map(I => gl_ram_n_58, ZN => CTS_297);
  CTS_ccl_a_BUF_clk_G0_L6_2 : CKBD2BWP7T port map(I => CTS_295, Z => CTS_294);
  CTS_cex_INV_clk_G0_L6_1 : CKND2BWP7T port map(I => CTS_295, ZN => CTS_293);
  CTS_ccl_a_BUF_clk_G0_L5_3 : CKBD6BWP7T port map(I => CTS_296, Z => CTS_295);
  CTS_cid_BUF_clk_G0_L4_4 : CKBD2BWP7T port map(I => gl_ram_n_56, Z => CTS_296);
  CTS_ccl_a_BUF_clk_G0_L5_2 : CKBD0BWP7T port map(I => CTS_292, Z => CTS_291);
  CTS_cex_INV_clk_G0_L5_1 : CKND0BWP7T port map(I => CTS_292, ZN => CTS_290);
  CTS_cid_BUF_clk_G0_L4_3 : CKBD2BWP7T port map(I => gl_ram_n_52, Z => CTS_292);
  CTS_ccl_a_BUF_clk_G0_L2_2 : CKBD12BWP7T port map(I => CTS_365, Z => CTS_345);
  CTS_ccl_a_BUF_clk_G0_L3_2 : CKBD8BWP7T port map(I => CTS_289, Z => CTS_288);
  CTS_ccl_a_BUF_clk_G0_L2_1 : CKBD6BWP7T port map(I => CTS_365, Z => CTS_289);
  CTS_ccl_a_BUF_clk_G0_L4_2 : CKBD0BWP7T port map(I => CTS_287, Z => CTS_286);
  CTS_cex_INV_clk_G0_L4_1 : CKND1BWP7T port map(I => CTS_287, ZN => CTS_285);
  CTS_ccl_a_BUF_clk_G0_L3_1 : CKBD0BWP7T port map(I => gl_ram_n_62, Z => CTS_287);
  CTS_ccl_a_BUF_clk_G0_L1_1 : CKBD4BWP7T port map(I => clk, Z => CTS_365);
  FE_OCPC159_gl_ram_ram_59_2 : BUFFD1BWP7T port map(I => gl_ram_ram_59(2), Z => FE_OCPN159_gl_ram_ram_59_2);
  FE_RC_74_0 : CKND2D3BWP7T port map(A1 => gl_ram_ram_81(0), A2 => gl_ram_n_88, ZN => FE_RN_23_0);
  FE_RC_73_0 : ND2D3BWP7T port map(A1 => FE_RN_23_0, A2 => gl_ram_n_251, ZN => gl_ram_n_1499);
  FE_RC_70_0 : AOI21D2BWP7T port map(A1 => gl_ram_n_1439, A2 => gl_ram_n_590, B => gl_ram_n_554, ZN => gl_ram_n_668);
  FE_RC_69_0 : ND2D2BWP7T port map(A1 => gl_ram_ram_88(2), A2 => gl_ram_n_89, ZN => FE_RN_21_0);
  FE_RC_68_0 : ND2D2BWP7T port map(A1 => gl_ram_n_336, A2 => FE_RN_21_0, ZN => gl_ram_n_1476);
  FE_RC_67_0 : ND2D2BWP7T port map(A1 => gl_ram_ram_16(2), A2 => gl_ram_n_89, ZN => FE_RN_20_0);
  FE_RC_66_0 : ND2D2BWP7T port map(A1 => FE_RN_20_0, A2 => gl_ram_n_311, ZN => gl_ram_n_1452);
  FE_RC_65_0 : ND2D2BWP7T port map(A1 => gl_ram_ram_70(2), A2 => gl_ram_n_93, ZN => FE_RN_19_0);
  FE_RC_64_0 : ND2D2BWP7T port map(A1 => FE_RN_19_0, A2 => gl_ram_n_357, ZN => gl_ram_n_1467);
  FE_RC_63_0 : INVD1BWP7T port map(I => gl_ram_n_86, ZN => FE_RN_18_0);
  FE_RC_62_0 : IND2D2BWP7T port map(A1 => FE_RN_18_0, B1 => gl_ram_ram_50(2), ZN => gl_ram_n_282);
  FE_RC_61_0 : INVD1BWP7T port map(I => gl_ram_n_90, ZN => FE_RN_16_0);
  FE_RC_60_0 : IND2D2BWP7T port map(A1 => FE_RN_16_0, B1 => gl_ram_ram_77(2), ZN => FE_RN_17_0);
  FE_RC_59_0 : ND2D2BWP7T port map(A1 => gl_ram_n_366, A2 => FE_RN_17_0, ZN => gl_ram_n_1463);
  FE_RC_58_0 : INVD1BWP7T port map(I => gl_ram_n_88, ZN => FE_RN_15_0);
  FE_RC_57_0 : IND2D2BWP7T port map(A1 => FE_RN_15_0, B1 => gl_ram_ram_49(2), ZN => gl_ram_n_281);
  FE_RC_56_0 : INVD1BWP7T port map(I => gl_ram_n_91, ZN => FE_RN_14_0);
  FE_RC_55_0 : IND2D2BWP7T port map(A1 => FE_RN_14_0, B1 => gl_ram_ram_52(2), ZN => gl_ram_n_283);
  FE_RC_54_0 : INVD1BWP7T port map(I => gl_ram_n_90, ZN => FE_RN_13_0);
  FE_OCPC151_gl_ram_ram_15_1 : BUFFD1BWP7T port map(I => gl_ram_ram_15(1), Z => FE_OCPN151_gl_ram_ram_15_1);
  FE_OCPC150_gl_ram_ram_23_1 : BUFFD1BWP7T port map(I => gl_ram_ram_23(1), Z => FE_OCPN150_gl_ram_ram_23_1);
  FE_RC_52_0 : INVD1BWP7T port map(I => gl_ram_n_555, ZN => FE_RN_11_0);
  FE_RC_51_0 : IND2D4BWP7T port map(A1 => FE_RN_11_0, B1 => gl_ram_n_657, ZN => FE_RN_12_0);
  FE_RC_50_0 : ND2D5BWP7T port map(A1 => FE_RN_12_0, A2 => gl_ram_n_7, ZN => gl_ram_n_699);
  FE_RC_49_0 : AOI21D2BWP7T port map(A1 => gl_ram_n_628, A2 => gl_ram_n_629, B => gl_ram_n_94, ZN => gl_ram_n_680);
  FE_RC_47_0 : ND2D2BWP7T port map(A1 => gl_ram_ram_89(2), A2 => gl_ram_n_88, ZN => FE_RN_10_0);
  FE_RC_46_0 : ND2D2BWP7T port map(A1 => gl_ram_n_339, A2 => FE_RN_10_0, ZN => gl_ram_n_1475);
  FE_RC_44_0 : CKND1BWP7T port map(I => gl_ram_n_561, ZN => FE_RN_8_0);
  FE_RC_43_0 : ND2D2BWP7T port map(A1 => gl_ram_n_592, A2 => gl_ram_n_593, ZN => FE_RN_9_0);
  FE_RC_42_0 : CKND2D3BWP7T port map(A1 => FE_RN_9_0, A2 => FE_RN_8_0, ZN => gl_ram_n_7);
  FE_OCPC148_gl_ram_ram_4_1 : BUFFD1BWP7T port map(I => gl_ram_ram_4(1), Z => FE_OCPN148_gl_ram_ram_4_1);
  FE_OCPC147_gl_ram_ram_6_1 : BUFFD1BWP7T port map(I => gl_ram_ram_6(1), Z => FE_OCPN147_gl_ram_ram_6_1);
  FE_OCPC146_gl_ram_ram_86_1 : BUFFD1BWP7T port map(I => gl_ram_ram_86(1), Z => FE_OCPN146_gl_ram_ram_86_1);
  FE_OCPC145_gl_ram_ram_88_1 : BUFFD0BWP7T port map(I => gl_ram_ram_88(1), Z => FE_OCPN145_gl_ram_ram_88_1);
  FE_OCPC144_gl_ram_ram_87_1 : BUFFD0BWP7T port map(I => gl_ram_ram_87(1), Z => FE_OCPN144_gl_ram_ram_87_1);
  FE_OCPC143_gl_ram_ram_3_1 : BUFFD1BWP7T port map(I => gl_ram_ram_3(1), Z => FE_OCPN143_gl_ram_ram_3_1);
  FE_OCPC140_gl_ram_ram_89_1 : BUFFD0BWP7T port map(I => gl_ram_ram_89(1), Z => FE_OCPN140_gl_ram_ram_89_1);
  FE_OCPC139_gl_ram_ram_90_1 : BUFFD0BWP7T port map(I => gl_ram_ram_90(1), Z => FE_OCPN139_gl_ram_ram_90_1);
  FE_OCPC136_gl_ram_ram_51_1 : BUFFD0BWP7T port map(I => gl_ram_ram_51(1), Z => FE_OCPN136_gl_ram_ram_51_1);
  FE_OCPC133_gl_ram_ram_76_1 : BUFFD0BWP7T port map(I => gl_ram_ram_76(1), Z => FE_OCPN133_gl_ram_ram_76_1);
  FE_OCPC130_gl_ram_ram_80_1 : BUFFD1BWP7T port map(I => gl_ram_ram_80(1), Z => FE_OCPN130_gl_ram_ram_80_1);
  FE_OCPC127_gl_ram_ram_81_1 : BUFFD1BWP7T port map(I => gl_ram_ram_81(1), Z => FE_OCPN127_gl_ram_ram_81_1);
  FE_OCPC126_gl_ram_ram_21_1 : BUFFD0BWP7T port map(I => gl_ram_ram_21(1), Z => FE_OCPN126_gl_ram_ram_21_1);
  FE_OCPC125_gl_ram_ram_67_1 : BUFFD0BWP7T port map(I => gl_ram_ram_67(1), Z => FE_OCPN125_gl_ram_ram_67_1);
  FE_OCPC123_gl_ram_ram_85_1 : BUFFD1BWP7T port map(I => gl_ram_ram_85(1), Z => FE_OCPN123_gl_ram_ram_85_1);
  FE_OCPC119_gl_ram_ram_91_1 : BUFFD0BWP7T port map(I => gl_ram_ram_91(1), Z => FE_OCPN119_gl_ram_ram_91_1);
  FE_OCPC117_gl_ram_ram_92_1 : BUFFD1BWP7T port map(I => gl_ram_ram_92(1), Z => FE_OCPN117_gl_ram_ram_92_1);
  FE_OCPC116_gl_ram_ram_71_1 : BUFFD1BWP7T port map(I => gl_ram_ram_71(1), Z => FE_OCPN116_gl_ram_ram_71_1);
  FE_OCPC111_gl_ram_ram_10_2 : BUFFD1BWP7T port map(I => gl_ram_ram_10(2), Z => FE_OCPN111_gl_ram_ram_10_2);
  FE_OCPC110_gl_ram_ram_77_1 : BUFFD0BWP7T port map(I => gl_ram_ram_77(1), Z => FE_OCPN110_gl_ram_ram_77_1);
  FE_OCPC108_gl_ram_ram_76_2 : BUFFD0BWP7T port map(I => gl_ram_ram_76(2), Z => FE_OCPN108_gl_ram_ram_76_2);
  FE_OCPC107_gl_ram_ram_78_1 : BUFFD1BWP7T port map(I => gl_ram_ram_78(1), Z => FE_OCPN107_gl_ram_ram_78_1);
  FE_OCPC103_gl_ram_ram_13_2 : BUFFD1BWP7T port map(I => FE_OCPN273_gl_ram_ram_13_2, Z => FE_OCPN103_gl_ram_ram_13_2);
  FE_OCPC102_gl_ram_ram_79_1 : BUFFD0BWP7T port map(I => gl_ram_ram_79(1), Z => FE_OCPN102_gl_ram_ram_79_1);
  FE_RC_39_0 : CKND2D2BWP7T port map(A1 => gl_ram_ram_13(1), A2 => gl_ram_n_90, ZN => FE_RN_7_0);
  FE_RC_38_0 : ND2D3BWP7T port map(A1 => FE_RN_7_0, A2 => gl_ram_n_401, ZN => gl_ram_n_1453);
  FE_OCPC89_gl_ram_ram_24_0 : BUFFD1BWP7T port map(I => gl_ram_ram_24(0), Z => FE_OCPN89_gl_ram_ram_24_0);
  FE_OCPC85_gl_ram_ram_14_2 : BUFFD1BWP7T port map(I => gl_ram_ram_14(2), Z => FE_OCPN85_gl_ram_ram_14_2);
  FE_OCPC77_gl_ram_ram_32_2 : BUFFD0BWP7T port map(I => gl_ram_ram_32(2), Z => FE_OCPN77_gl_ram_ram_32_2);
  FE_OCPC74_gl_ram_ram_21_0 : BUFFD1BWP7T port map(I => gl_ram_ram_21(0), Z => FE_OCPN74_gl_ram_ram_21_0);
  FE_RC_37_0 : IOA21D2BWP7T port map(A1 => gl_ram_ram_59(2), A2 => gl_ram_n_87, B => FE_RN_5_0, ZN => gl_ram_n_1478);
  FE_OCPC72_gl_ram_ram_8_1 : BUFFD1BWP7T port map(I => gl_ram_ram_8(1), Z => FE_OCPN72_gl_ram_ram_8_1);
  FE_OCPC71_gl_ram_ram_1_1 : BUFFD1BWP7T port map(I => gl_ram_ram_1(1), Z => FE_OCPN71_gl_ram_ram_1_1);
  FE_OCPC70_gl_ram_ram_73_1 : BUFFD0BWP7T port map(I => gl_ram_ram_73(1), Z => FE_OCPN70_gl_ram_ram_73_1);
  FE_OCPC67_gl_ram_ram_77_0 : BUFFD1BWP7T port map(I => gl_ram_ram_77(0), Z => FE_OCPN67_gl_ram_ram_77_0);
  FE_RC_35_0 : ND2D2BWP7T port map(A1 => gl_ram_ram_57(1), A2 => gl_ram_n_88, ZN => FE_RN_6_0);
  FE_RC_34_0 : IOA21D2BWP7T port map(A1 => gl_ram_ram_58(1), A2 => gl_ram_n_86, B => FE_RN_6_0, ZN => gl_ram_n_426);
  FE_OCPC66_gl_ram_ram_29_0 : BUFFD0BWP7T port map(I => gl_ram_ram_29(0), Z => FE_OCPN66_gl_ram_ram_29_0);
  FE_OCPC65_gl_ram_ram_74_1 : BUFFD1BWP7T port map(I => gl_ram_ram_74(1), Z => FE_OCPN65_gl_ram_ram_74_1);
  FE_OCPC63_gl_ram_ram_31_0 : BUFFD1BWP7T port map(I => gl_ram_ram_31(0), Z => FE_OCPN63_gl_ram_ram_31_0);
  FE_OCPC61_gl_ram_ram_55_2 : BUFFD1BWP7T port map(I => FE_PSN350_gl_ram_ram_55_2, Z => FE_OCPN61_gl_ram_ram_55_2);
  FE_OCPC56_gl_ram_ram_33_1 : BUFFD0BWP7T port map(I => gl_ram_ram_33(1), Z => FE_OCPN56_gl_ram_ram_33_1);
  FE_OCPC54_gl_ram_ram_48_1 : BUFFD1BWP7T port map(I => gl_ram_ram_48(1), Z => FE_OCPN54_gl_ram_ram_48_1);
  FE_OCPC46_gl_ram_ram_41_0 : BUFFD1BWP7T port map(I => gl_ram_ram_41(0), Z => FE_OCPN46_gl_ram_ram_41_0);
  FE_OCPC43_gl_ram_ram_56_0 : BUFFD1BWP7T port map(I => gl_ram_ram_56(0), Z => FE_OCPN43_gl_ram_ram_56_0);
  FE_OCPC42_gl_ram_ram_60_0 : BUFFD1BWP7T port map(I => gl_ram_ram_60(0), Z => FE_OCPN42_gl_ram_ram_60_0);
  FE_OCPC38_gl_ram_ram_48_0 : BUFFD0BWP7T port map(I => gl_ram_ram_48(0), Z => FE_OCPN38_gl_ram_ram_48_0);
  FE_OCPC28_gl_ram_ram_10_1 : BUFFD0BWP7T port map(I => gl_ram_ram_10(1), Z => FE_OCPN28_gl_ram_ram_10_1);
  FE_OCPC14_gl_ram_ram_28_1 : BUFFD1BWP7T port map(I => gl_ram_ram_28(1), Z => FE_OCPN14_gl_ram_ram_28_1);
  FE_OCPC10_gl_ram_ram_25_1 : BUFFD0BWP7T port map(I => gl_ram_ram_25(1), Z => FE_OCPN10_gl_ram_ram_25_1);
  FE_OCPC8_gl_ram_ram_47_1 : BUFFD1BWP7T port map(I => gl_ram_ram_47(1), Z => FE_OCPN8_gl_ram_ram_47_1);
  FE_RC_31_0 : ND2D2BWP7T port map(A1 => gl_ram_ram_56(2), A2 => gl_ram_n_89, ZN => FE_RN_5_0);
  FE_OCPC7_gl_ram_ram_40_1 : BUFFD0BWP7T port map(I => gl_ram_ram_40(1), Z => FE_OCPN7_gl_ram_ram_40_1);
  FE_OCPC6_gl_ram_ram_30_1 : BUFFD1BWP7T port map(I => gl_ram_ram_30(1), Z => FE_OCPN6_gl_ram_ram_30_1);
  FE_RC_29_0 : AOI21D2BWP7T port map(A1 => gl_ram_n_601, A2 => gl_ram_n_600, B => gl_ram_n_96, ZN => gl_ram_n_681);
  FE_OCPC2_gl_ram_ram_41_1 : BUFFD1BWP7T port map(I => gl_ram_ram_41(1), Z => FE_OCPN2_gl_ram_ram_41_1);
  FE_RC_25_0 : AOI21D2BWP7T port map(A1 => gl_ram_n_580, A2 => gl_ram_n_579, B => gl_ram_n_94, ZN => gl_ram_n_678);
  FE_RC_24_0 : AOI21D2BWP7T port map(A1 => gl_ram_n_607, A2 => gl_ram_n_606, B => gl_ram_n_107, ZN => gl_ram_n_691);
  FE_RC_20_0 : AOI21D2BWP7T port map(A1 => gl_ram_n_645, A2 => gl_ram_n_644, B => gl_ram_n_98, ZN => gl_ram_n_677);
  FE_RC_19_0 : AOI21D2BWP7T port map(A1 => gl_ram_n_623, A2 => gl_ram_n_624, B => gl_ram_n_99, ZN => gl_ram_n_687);
  FE_RC_17_0 : ND2D3BWP7T port map(A1 => gl_ram_n_639, A2 => gl_ram_n_638, ZN => FE_RN_3_0);
  FE_RC_16_0 : CKND2D4BWP7T port map(A1 => FE_RN_3_0, A2 => gl_ram_n_559, ZN => gl_ram_n_1549);
  FE_OCPC3_gl_ram_n_1448 : INVD6BWP7T port map(I => FE_OCPN0_gl_ram_n_1448, ZN => FE_OCPN3_gl_ram_n_1448);
  FE_OCPC2_gl_ram_n_1448 : INVD6BWP7T port map(I => FE_OCPN0_gl_ram_n_1448, ZN => FE_OCPN2_gl_ram_n_1448);
  FE_OCPC1_gl_ram_n_1448 : INVD4BWP7T port map(I => FE_OCPN0_gl_ram_n_1448, ZN => FE_OCPN1_gl_ram_n_1448);
  FE_OCPC0_gl_ram_n_1448 : CKND10BWP7T port map(I => gl_ram_n_1448, ZN => FE_OCPN0_gl_ram_n_1448);
  FE_RC_15_0 : AOI21D2BWP7T port map(A1 => gl_ram_n_626, A2 => gl_ram_n_627, B => gl_ram_n_96, ZN => gl_ram_n_682);
  FE_RC_14_0 : AOI21D2BWP7T port map(A1 => gl_ram_n_632, A2 => gl_ram_n_633, B => gl_ram_n_107, ZN => gl_ram_n_692);
  FE_RC_13_0 : CKND1BWP7T port map(I => gl_ram_n_560, ZN => FE_RN_1_0);
  FE_RC_12_0 : ND2D4BWP7T port map(A1 => gl_ram_n_641, A2 => gl_ram_n_640, ZN => FE_RN_2_0);
  FE_RC_11_0 : CKND2D4BWP7T port map(A1 => FE_RN_2_0, A2 => FE_RN_1_0, ZN => gl_ram_n_11);
  FE_RC_8_0 : AOI21D2BWP7T port map(A1 => gl_ram_n_587, A2 => gl_ram_n_588, B => gl_ram_n_552, ZN => gl_ram_n_665);
  FE_RC_7_0 : AOI21D2BWP7T port map(A1 => gl_ram_n_636, A2 => gl_ram_n_637, B => gl_ram_n_558, ZN => gl_ram_n_669);
  FE_RC_6_0 : ND2D1P5BWP7T port map(A1 => gl_ram_n_610, A2 => gl_ram_n_589, ZN => FE_RN_0_0);
  FE_RC_5_0 : CKND2D2BWP7T port map(A1 => FE_RN_0_0, A2 => gl_ram_n_553, ZN => gl_ram_n_1550);
  FE_RC_4_0 : ND4D4BWP7T port map(A1 => gl_ram_n_713, A2 => gl_ram_n_703, A3 => gl_ram_n_704, A4 => gl_ram_n_702, ZN => gl_ram_n_720);
  FE_RC_3_0 : AOI21D2BWP7T port map(A1 => gl_ram_n_620, A2 => gl_ram_n_621, B => gl_ram_n_4, ZN => gl_ram_n_694);
  FE_RC_1_0 : AOI21D2BWP7T port map(A1 => gl_ram_n_575, A2 => gl_ram_n_659, B => gl_ram_n_408, ZN => gl_ram_n_708);
  FE_DBTC0_reset : INVD1P5BWP7T port map(I => FE_OFN31_reset, ZN => FE_DBTN0_reset);
  gl_g1475 : ND3D0BWP7T port map(A1 => gl_n_45, A2 => gl_n_36, A3 => gl_n_42, ZN => gl_sig_green);
  gl_g1476 : IND4D0BWP7T port map(A1 => gl_sig_y(2), B1 => gl_sig_y(1), B2 => gl_sig_y(0), B3 => gl_n_44, ZN => gl_n_45);
  gl_g1477 : NR4D0BWP7T port map(A1 => gl_n_31, A2 => gl_n_43, A3 => gl_n_24, A4 => gl_sig_y(3), ZN => gl_n_44);
  gl_g1478 : OAI221D0BWP7T port map(A1 => gl_n_39, A2 => gl_n_38, B1 => gl_n_27, B2 => gl_gr_lg_sig_countdown_5_141, C => gl_n_34, ZN => gl_n_43);
  gl_g1479 : CKND2D1BWP7T port map(A1 => gl_n_36, A2 => gl_n_41, ZN => gl_sig_blue);
  gl_g1480 : CKND2D1BWP7T port map(A1 => gl_n_36, A2 => gl_n_40, ZN => gl_sig_red);
  gl_g1481 : AOI22D0BWP7T port map(A1 => gl_sig_ram(1), A2 => gl_n_37, B1 => gl_n_33, B2 => sig_output_color(1), ZN => gl_n_42);
  gl_g1482 : AOI22D0BWP7T port map(A1 => gl_sig_ram(2), A2 => gl_n_37, B1 => gl_n_33, B2 => sig_output_color(2), ZN => gl_n_41);
  gl_g1483 : AOI22D0BWP7T port map(A1 => gl_sig_ram(0), A2 => gl_n_37, B1 => gl_n_33, B2 => sig_output_color(0), ZN => gl_n_40);
  gl_g1484 : OAI32D1BWP7T port map(A1 => gl_n_32, A2 => gl_n_28, A3 => gl_n_25, B1 => gl_n_29, B2 => gl_n_4, ZN => gl_n_39);
  gl_g1485 : NR3D0BWP7T port map(A1 => gl_n_32, A2 => gl_n_3, A3 => gl_n_22, ZN => gl_n_38);
  gl_g1486 : AOI211XD0BWP7T port map(A1 => gl_n_19, A2 => gl_sig_x(3), B => gl_n_35, C => gl_n_21, ZN => gl_n_37);
  gl_g1487 : ND2D1BWP7T port map(A1 => gl_n_33, A2 => gl_sig_rom(0), ZN => gl_n_36);
  gl_g1488 : OAI22D0BWP7T port map(A1 => gl_sig_rom(0), A2 => gl_n_30, B1 => gl_n_16, B2 => gl_sig_y(3), ZN => gl_n_35);
  gl_g1489 : AOI22D0BWP7T port map(A1 => gl_gr_lg_sig_countdown_7_139, A2 => gl_n_27, B1 => gl_gr_lg_sig_countdown_5_141, B2 => gl_n_2, ZN => gl_n_34);
  gl_g1490 : INR2D1BWP7T port map(A1 => gl_sig_rom(1), B1 => gl_n_30, ZN => gl_n_33);
  gl_g1491 : NR2D0BWP7T port map(A1 => gl_sig_rom(0), A2 => gl_n_30, ZN => gl_n_31);
  gl_g1492 : INR2D0BWP7T port map(A1 => gl_n_29, B1 => gl_sig_x(3), ZN => gl_n_32);
  gl_g1493 : ND4D0BWP7T port map(A1 => gl_n_26, A2 => gl_n_14, A3 => gl_n_12, A4 => gl_gr_lg_le_n_22, ZN => gl_n_30);
  gl_g1494 : OAI21D0BWP7T port map(A1 => gl_gr_lg_sig_countdown_4_142, A2 => gl_n_20, B => gl_n_27, ZN => gl_n_29);
  gl_g1495 : MOAI22D0BWP7T port map(A1 => gl_sig_x(0), A2 => gl_n_6, B1 => gl_n_3, B2 => gl_n_22, ZN => gl_n_28);
  gl_g1496 : ND2D0BWP7T port map(A1 => gl_gr_lg_sig_countdown_4_142, A2 => gl_n_20, ZN => gl_n_27);
  gl_g1497 : NR4D0BWP7T port map(A1 => gl_n_23, A2 => gl_n_8, A3 => gl_n_9, A4 => gl_n_10, ZN => gl_n_26);
  gl_g1498 : AOI21D0BWP7T port map(A1 => gl_n_15, A2 => gl_n_6, B => gl_sig_x(1), ZN => gl_n_25);
  gl_g1499 : OAI22D0BWP7T port map(A1 => gl_n_18, A2 => gl_sig_x(0), B1 => gl_n_2, B2 => gl_gr_lg_sig_countdown_7_139, ZN => gl_n_24);
  gl_g1500 : OAI211D1BWP7T port map(A1 => sig_logic_x(1), A2 => gl_n_0, B => gl_n_11, C => gl_n_7, ZN => gl_n_23);
  gl_g1501 : NR4D0BWP7T port map(A1 => gl_sig_x(1), A2 => gl_sig_x(2), A3 => gl_sig_x(0), A4 => gl_sig_x(3), ZN => gl_n_21);
  gl_g1502 : AO21D0BWP7T port map(A1 => gl_n_1, A2 => gl_n_6, B => gl_n_20, Z => gl_n_22);
  gl_g1503 : IOA21D1BWP7T port map(A1 => gl_sig_x(1), A2 => gl_sig_x(0), B => gl_n_3, ZN => gl_n_19);
  gl_g1504 : ND3D0BWP7T port map(A1 => gl_sig_x(1), A2 => gl_sig_x(3), A3 => gl_sig_x(2), ZN => gl_n_18);
  gl_g1505 : OA21D0BWP7T port map(A1 => gl_sig_y(1), A2 => gl_sig_y(0), B => gl_sig_y(2), Z => gl_n_16);
  gl_g1506 : MAOI22D0BWP7T port map(A1 => gl_n_5, A2 => gl_gr_lg_sig_countdown_1_145, B1 => gl_gr_lg_sig_countdown_2_144, B2 => gl_gr_lg_sig_countdown_1_145, ZN => gl_n_15);
  gl_g1507 : XNR2D1BWP7T port map(A1 => sig_logic_y(1), A2 => gl_sig_y(1), ZN => gl_n_14);
  gl_g1508 : NR2D0BWP7T port map(A1 => gl_n_1, A2 => gl_n_6, ZN => gl_n_20);
  gl_g1510 : XNR2D1BWP7T port map(A1 => sig_logic_y(0), A2 => gl_sig_y(0), ZN => gl_n_12);
  gl_g1511 : XNR2D1BWP7T port map(A1 => sig_logic_y(3), A2 => gl_sig_y(3), ZN => gl_n_11);
  gl_g1512 : MOAI22D0BWP7T port map(A1 => gl_n_5, A2 => sig_logic_x(0), B1 => gl_n_5, B2 => FE_PHN505_sig_logic_x_0, ZN => gl_n_10);
  gl_g1513 : MOAI22D0BWP7T port map(A1 => gl_n_4, A2 => sig_logic_x(3), B1 => gl_n_4, B2 => sig_logic_x(3), ZN => gl_n_9);
  gl_g1514 : MOAI22D0BWP7T port map(A1 => gl_n_3, A2 => sig_logic_x(2), B1 => gl_n_3, B2 => sig_logic_x(2), ZN => gl_n_8);
  gl_g1515 : CKND2D0BWP7T port map(A1 => gl_n_0, A2 => sig_logic_x(1), ZN => gl_n_7);
  gl_g1516 : ND2D0BWP7T port map(A1 => gl_gr_lg_sig_countdown_2_144, A2 => gl_gr_lg_sig_countdown_1_145, ZN => gl_n_6);
  gl_g1517 : INVD1BWP7T port map(I => gl_sig_x(0), ZN => gl_n_5);
  gl_g1518 : INVD1BWP7T port map(I => gl_sig_x(3), ZN => gl_n_4);
  gl_g1519 : INVD1BWP7T port map(I => gl_sig_x(2), ZN => gl_n_3);
  gl_g1520 : CKND1BWP7T port map(I => gl_gr_lg_sig_countdown_6_140, ZN => gl_n_2);
  gl_g1521 : CKND1BWP7T port map(I => gl_gr_lg_sig_countdown_3_143, ZN => gl_n_1);
  gl_g1522 : INVD1BWP7T port map(I => gl_sig_x(1), ZN => gl_n_0);
  gl_gr_lg_le_g55 : INVD0BWP7T port map(I => gl_gr_lg_le_n_32, ZN => gl_gr_lg_le_n_31);
  gl_gr_lg_le_g270 : AN4D1BWP7T port map(A1 => gl_gr_lg_le_n_29, A2 => gl_gr_lg_le_n_24, A3 => gl_gr_lg_le_n_25, A4 => gl_gr_lg_le_n_20, Z => gl_gr_lg_le_n_32);
  gl_gr_lg_le_g271 : NR4D0BWP7T port map(A1 => gl_gr_lg_le_n_28, A2 => gl_gr_lg_le_n_26, A3 => gl_gr_lg_le_n_23, A4 => gl_gr_lg_le_n_21, ZN => gl_gr_lg_le_n_29);
  gl_gr_lg_le_g272 : ND2D1BWP7T port map(A1 => gl_gr_lg_le_n_27, A2 => gl_gr_lg_le_n_22, ZN => gl_gr_lg_le_n_28);
  gl_gr_lg_le_g273 : XNR2D1BWP7T port map(A1 => sig_logic_x(2), A2 => gl_sig_x(2), ZN => gl_gr_lg_le_n_27);
  gl_gr_lg_le_g274 : CKXOR2D0BWP7T port map(A1 => sig_logic_x(3), A2 => gl_sig_x(3), Z => gl_gr_lg_le_n_26);
  gl_gr_lg_le_g275 : MOAI22D0BWP7T port map(A1 => sig_logic_y(0), A2 => gl_sig_y(0), B1 => sig_logic_y(0), B2 => gl_sig_y(0), ZN => gl_gr_lg_le_n_25);
  gl_gr_lg_le_g276 : MOAI22D0BWP7T port map(A1 => FE_PHN316_sig_logic_y_3, A2 => gl_sig_y(3), B1 => FE_PHN316_sig_logic_y_3, B2 => gl_sig_y(3), ZN => gl_gr_lg_le_n_24);
  gl_gr_lg_le_g277 : CKXOR2D0BWP7T port map(A1 => sig_logic_x(0), A2 => gl_sig_x(0), Z => gl_gr_lg_le_n_23);
  gl_gr_lg_le_g278 : XNR2D1BWP7T port map(A1 => sig_logic_y(2), A2 => gl_sig_y(2), ZN => gl_gr_lg_le_n_22);
  gl_gr_lg_le_g279 : CKXOR2D0BWP7T port map(A1 => sig_logic_x(1), A2 => gl_sig_x(1), Z => gl_gr_lg_le_n_21);
  gl_gr_lg_le_g280 : MOAI22D0BWP7T port map(A1 => sig_logic_y(1), A2 => gl_sig_y(1), B1 => sig_logic_y(1), B2 => gl_sig_y(1), ZN => gl_gr_lg_le_n_20);
  gl_gr_lg_le_new_count_e_reg_9 : LNQD1BWP7T port map(D => gl_gr_lg_le_n_19, EN => gl_gr_lg_le_n_18, Q => gl_gr_lg_le_new_count_e(9));
  gl_gr_lg_le_g292 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_le_n_16, A2 => gl_sig_e(9), B1 => gl_gr_lg_le_n_16, B2 => gl_sig_e(9), ZN => gl_gr_lg_le_n_19);
  gl_gr_lg_le_new_count_e_reg_8 : LNQD1BWP7T port map(D => gl_gr_lg_le_n_17, EN => gl_gr_lg_le_n_18, Q => gl_gr_lg_le_new_count_e(8));
  gl_gr_lg_le_g294 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_le_n_14, A2 => gl_sig_e(8), B1 => gl_gr_lg_le_n_14, B2 => gl_sig_e(8), ZN => gl_gr_lg_le_n_17);
  gl_gr_lg_le_new_count_e_reg_7 : LNQD1BWP7T port map(D => gl_gr_lg_le_n_15, EN => gl_gr_lg_le_n_18, Q => gl_gr_lg_le_new_count_e(7));
  gl_gr_lg_le_g296 : IND2D1BWP7T port map(A1 => gl_gr_lg_le_n_14, B1 => gl_sig_e(8), ZN => gl_gr_lg_le_n_16);
  gl_gr_lg_le_g297 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_le_n_12, A2 => gl_sig_e(7), B1 => gl_gr_lg_le_n_12, B2 => gl_sig_e(7), ZN => gl_gr_lg_le_n_15);
  gl_gr_lg_le_new_count_e_reg_6 : LNQD1BWP7T port map(D => gl_gr_lg_le_n_13, EN => gl_gr_lg_le_n_18, Q => gl_gr_lg_le_new_count_e(6));
  gl_gr_lg_le_g299 : IND2D1BWP7T port map(A1 => gl_gr_lg_le_n_12, B1 => gl_sig_e(7), ZN => gl_gr_lg_le_n_14);
  gl_gr_lg_le_g300 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_le_n_10, A2 => gl_sig_e(6), B1 => gl_gr_lg_le_n_10, B2 => gl_sig_e(6), ZN => gl_gr_lg_le_n_13);
  gl_gr_lg_le_new_count_e_reg_5 : LNQD1BWP7T port map(D => gl_gr_lg_le_n_11, EN => gl_gr_lg_le_n_18, Q => gl_gr_lg_le_new_count_e(5));
  gl_gr_lg_le_g302 : IND2D1BWP7T port map(A1 => gl_gr_lg_le_n_10, B1 => gl_sig_e(6), ZN => gl_gr_lg_le_n_12);
  gl_gr_lg_le_g303 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_le_n_8, A2 => gl_sig_e(5), B1 => gl_gr_lg_le_n_8, B2 => gl_sig_e(5), ZN => gl_gr_lg_le_n_11);
  gl_gr_lg_le_new_count_e_reg_4 : LNQD1BWP7T port map(D => gl_gr_lg_le_n_9, EN => gl_gr_lg_le_n_18, Q => gl_gr_lg_le_new_count_e(4));
  gl_gr_lg_le_g305 : IND2D1BWP7T port map(A1 => gl_gr_lg_le_n_8, B1 => gl_sig_e(5), ZN => gl_gr_lg_le_n_10);
  gl_gr_lg_le_g306 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_le_n_6, A2 => gl_sig_e(4), B1 => gl_gr_lg_le_n_6, B2 => gl_sig_e(4), ZN => gl_gr_lg_le_n_9);
  gl_gr_lg_le_new_count_e_reg_3 : LNQD1BWP7T port map(D => gl_gr_lg_le_n_7, EN => gl_gr_lg_le_n_18, Q => gl_gr_lg_le_new_count_e(3));
  gl_gr_lg_le_g308 : IND2D1BWP7T port map(A1 => gl_gr_lg_le_n_6, B1 => gl_sig_e(4), ZN => gl_gr_lg_le_n_8);
  gl_gr_lg_le_g309 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_le_n_4, A2 => gl_sig_e(3), B1 => gl_gr_lg_le_n_4, B2 => gl_sig_e(3), ZN => gl_gr_lg_le_n_7);
  gl_gr_lg_le_new_count_e_reg_2 : LNQD1BWP7T port map(D => gl_gr_lg_le_n_5, EN => gl_gr_lg_le_n_18, Q => gl_gr_lg_le_new_count_e(2));
  gl_gr_lg_le_g311 : IND2D1BWP7T port map(A1 => gl_gr_lg_le_n_4, B1 => gl_sig_e(3), ZN => gl_gr_lg_le_n_6);
  gl_gr_lg_le_g312 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_le_n_2, A2 => gl_sig_e(2), B1 => gl_gr_lg_le_n_2, B2 => gl_sig_e(2), ZN => gl_gr_lg_le_n_5);
  gl_gr_lg_le_new_count_e_reg_1 : LNQD1BWP7T port map(D => gl_gr_lg_le_n_3, EN => gl_gr_lg_le_n_18, Q => FE_PHN376_gl_gr_lg_le_new_count_e_1);
  gl_gr_lg_le_g314 : IND2D1BWP7T port map(A1 => gl_gr_lg_le_n_2, B1 => gl_sig_e(2), ZN => gl_gr_lg_le_n_4);
  gl_gr_lg_le_g315 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_le_n_0, A2 => gl_sig_e(1), B1 => gl_gr_lg_le_n_0, B2 => gl_sig_e(1), ZN => gl_gr_lg_le_n_3);
  gl_gr_lg_le_new_count_e_reg_0 : LNQD1BWP7T port map(D => gl_gr_lg_le_n_1, EN => gl_gr_lg_le_n_18, Q => gl_gr_lg_le_new_count_e(0));
  gl_gr_lg_le_g317 : IND2D1BWP7T port map(A1 => gl_gr_lg_le_n_0, B1 => gl_sig_e(1), ZN => gl_gr_lg_le_n_2);
  gl_gr_lg_le_count_e_reg_9 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_322, D => FE_PHN372_gl_gr_lg_le_new_count_e_9, Q => gl_sig_e(9));
  gl_gr_lg_le_count_e_reg_5 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_322, D => FE_PHN369_gl_gr_lg_le_new_count_e_5, Q => gl_sig_e(5));
  gl_gr_lg_le_count_e_reg_6 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_322, D => FE_PHN374_gl_gr_lg_le_new_count_e_6, Q => gl_sig_e(6));
  gl_gr_lg_le_count_e_reg_8 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_322, D => FE_PHN373_gl_gr_lg_le_new_count_e_8, Q => gl_sig_e(8));
  gl_gr_lg_le_count_e_reg_7 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_322, D => FE_PHN371_gl_gr_lg_le_new_count_e_7, Q => gl_sig_e(7));
  gl_gr_lg_le_count_e_reg_1 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_322, D => gl_gr_lg_le_new_count_e(1), Q => gl_sig_e(1));
  gl_gr_lg_le_g324 : CKXOR2D1BWP7T port map(A1 => gl_gr_lg_le_n_32, A2 => gl_sig_e(0), Z => gl_gr_lg_le_n_1);
  gl_gr_lg_le_count_e_reg_2 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_322, D => FE_PHN363_gl_gr_lg_le_new_count_e_2, Q => gl_sig_e(2));
  gl_gr_lg_le_count_e_reg_3 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_322, D => FE_PHN366_gl_gr_lg_le_new_count_e_3, Q => gl_sig_e(3));
  gl_gr_lg_le_count_e_reg_4 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_322, D => FE_PHN364_gl_gr_lg_le_new_count_e_4, Q => gl_sig_e(4));
  gl_gr_lg_le_count_e_reg_0 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_322, D => FE_PHN367_gl_gr_lg_le_new_count_e_0, Q => gl_sig_e(0));
  gl_gr_lg_le_g329 : AOI21D2BWP7T port map(A1 => CTS_289, A2 => gl_gr_lg_le_n_32, B => gl_gr_lg_le_n_31, ZN => gl_gr_lg_le_n_18);
  gl_gr_lg_le_g330 : ND2D1BWP7T port map(A1 => gl_gr_lg_le_n_32, A2 => gl_sig_e(0), ZN => gl_gr_lg_le_n_0);
  gl_gr_lg_lv_g329 : OAI32D1BWP7T port map(A1 => gl_sig_y(2), A2 => gl_gr_lg_lv_n_3, A3 => gl_gr_lg_lv_n_7, B1 => gl_gr_lg_lv_n_1, B2 => gl_gr_lg_lv_n_12, ZN => gl_gr_lg_lv_n_14);
  gl_gr_lg_lv_g330 : OAI22D0BWP7T port map(A1 => gl_gr_lg_lv_n_12, A2 => gl_gr_lg_lv_n_2, B1 => gl_gr_lg_lv_n_7, B2 => gl_gr_lg_lv_n_9, ZN => FE_PHN400_gl_gr_lg_lv_n_13);
  gl_gr_lg_lv_count_v_reg_1 : DFQD1BWP7T port map(CP => CTS_288, D => FE_PHN426_gl_gr_lg_lv_n_10, Q => gl_sig_y(1));
  gl_gr_lg_lv_count_v_reg_0 : DFQD1BWP7T port map(CP => CTS_288, D => FE_PHN430_gl_gr_lg_lv_n_11, Q => gl_sig_y(0));
  gl_gr_lg_lv_g333 : AOI21D0BWP7T port map(A1 => gl_gr_lg_lv_n_6, A2 => gl_gr_lg_lv_n_3, B => gl_gr_lg_lv_n_8, ZN => gl_gr_lg_lv_n_12);
  gl_gr_lg_lv_g334 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_lv_n_7, A2 => gl_sig_y(0), B1 => gl_gr_lg_lv_n_8, B2 => gl_sig_y(0), ZN => gl_gr_lg_lv_n_11);
  gl_gr_lg_lv_g335 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_lv_n_7, A2 => gl_gr_lg_lv_n_0, B1 => gl_gr_lg_lv_n_8, B2 => gl_sig_y(1), ZN => gl_gr_lg_lv_n_10);
  gl_gr_lg_lv_g336 : OA32D1BWP7T port map(A1 => gl_sig_y(3), A2 => gl_gr_lg_lv_n_1, A3 => gl_gr_lg_lv_n_3, B1 => gl_sig_y(2), B2 => gl_gr_lg_lv_n_2, Z => gl_gr_lg_lv_n_9);
  gl_gr_lg_lv_g337 : NR2D1BWP7T port map(A1 => gl_gr_lg_lv_n_5, A2 => gl_gr_lg_lv_sig_edges, ZN => gl_gr_lg_lv_n_8);
  gl_gr_lg_lv_g338 : INVD1BWP7T port map(I => gl_gr_lg_lv_n_6, ZN => gl_gr_lg_lv_n_7);
  gl_gr_lg_lv_g339 : INR2XD0BWP7T port map(A1 => gl_gr_lg_lv_sig_edges, B1 => gl_gr_lg_lv_n_5, ZN => gl_gr_lg_lv_n_6);
  gl_gr_lg_lv_g340 : IND2D1BWP7T port map(A1 => FE_OFN31_reset, B1 => gl_gr_lg_lv_n_4, ZN => gl_gr_lg_lv_n_5);
  gl_gr_lg_lv_g341 : IND4D0BWP7T port map(A1 => gl_sig_y(0), B1 => gl_sig_y(3), B2 => gl_sig_y(2), B3 => gl_sig_y(1), ZN => gl_gr_lg_lv_n_4);
  gl_gr_lg_lv_g343 : ND2D1BWP7T port map(A1 => gl_sig_y(1), A2 => gl_sig_y(0), ZN => gl_gr_lg_lv_n_3);
  gl_gr_lg_lv_g2 : XNR2D1BWP7T port map(A1 => gl_sig_y(1), A2 => gl_sig_y(0), ZN => gl_gr_lg_lv_n_0);
  gl_gr_lg_lv_count_v_reg_3 : DFD1BWP7T port map(CP => CTS_288, D => gl_gr_lg_lv_n_13, Q => gl_sig_y(3), QN => gl_gr_lg_lv_n_2);
  gl_gr_lg_lv_count_v_reg_2 : DFD1BWP7T port map(CP => CTS_288, D => FE_PHN405_gl_gr_lg_lv_n_14, Q => gl_sig_y(2), QN => gl_gr_lg_lv_n_1);
  gl_gr_lg_lv_l_edge_g12 : NR2XD0BWP7T port map(A1 => gl_gr_lg_lv_l_edge_n_0, A2 => gl_gr_lg_lv_l_edge_reg2, ZN => gl_gr_lg_lv_sig_edges);
  gl_gr_lg_lv_l_edge_reg2_reg : DFQD1BWP7T port map(CP => CTS_288, D => FE_PHN368_gl_gr_lg_lv_l_edge_reg1, Q => gl_gr_lg_lv_l_edge_reg2);
  gl_gr_lg_lv_l_edge_reg1_reg : DFD1BWP7T port map(CP => CTS_288, D => FE_PHN382_gl_sig_scale_v, Q => gl_gr_lg_lv_l_edge_reg1, QN => gl_gr_lg_lv_l_edge_n_0);
  gl_gr_lg_lh_count_h_reg_3 : DFQD1BWP7T port map(CP => CTS_288, D => FE_PHN389_gl_gr_lg_lh_n_15, Q => gl_sig_x(3));
  gl_gr_lg_lh_g465 : OAI31D0BWP7T port map(A1 => gl_gr_lg_lh_n_2, A2 => gl_gr_lg_lh_n_0, A3 => gl_gr_lg_lh_n_5, B => gl_gr_lg_lh_n_12, ZN => gl_gr_lg_lh_n_15);
  gl_gr_lg_lh_g466 : OAI31D0BWP7T port map(A1 => gl_sig_x(2), A2 => gl_gr_lg_lh_n_2, A3 => gl_gr_lg_lh_n_5, B => gl_gr_lg_lh_n_13, ZN => gl_gr_lg_lh_n_14);
  gl_gr_lg_lh_g467 : ND2D1BWP7T port map(A1 => gl_gr_lg_lh_n_10, A2 => gl_sig_x(2), ZN => gl_gr_lg_lh_n_13);
  gl_gr_lg_lh_g468 : OAI21D0BWP7T port map(A1 => gl_gr_lg_lh_n_8, A2 => gl_gr_lg_lh_n_4, B => gl_sig_x(3), ZN => gl_gr_lg_lh_n_12);
  gl_gr_lg_lh_g469 : OAI22D0BWP7T port map(A1 => gl_gr_lg_lh_n_7, A2 => gl_gr_lg_lh_n_2, B1 => gl_gr_lg_lh_n_5, B2 => gl_sig_x(1), ZN => FE_PHN403_gl_gr_lg_lh_n_11);
  gl_gr_lg_lh_g471 : IOA21D1BWP7T port map(A1 => gl_gr_lg_lh_n_4, A2 => gl_gr_lg_lh_n_2, B => gl_gr_lg_lh_n_7, ZN => gl_gr_lg_lh_n_10);
  gl_gr_lg_lh_g472 : IOA21D1BWP7T port map(A1 => gl_sig_x(0), A2 => gl_gr_lg_lh_n_3, B => gl_gr_lg_lh_n_6, ZN => gl_gr_lg_lh_n_9);
  gl_gr_lg_lh_g473 : INVD1BWP7T port map(I => gl_gr_lg_lh_n_7, ZN => gl_gr_lg_lh_n_8);
  gl_gr_lg_lh_g474 : AOI21D0BWP7T port map(A1 => gl_gr_lg_lh_n_4, A2 => gl_gr_lg_lh_n_1, B => gl_gr_lg_lh_n_3, ZN => gl_gr_lg_lh_n_7);
  gl_gr_lg_lh_g475 : ND3D0BWP7T port map(A1 => gl_gr_lg_lh_n_4, A2 => gl_gr_lg_lh_n_1, A3 => gl_gr_lg_lh_sig_edges, ZN => gl_gr_lg_lh_n_6);
  gl_gr_lg_lh_g476 : ND3D0BWP7T port map(A1 => gl_gr_lg_lh_n_4, A2 => gl_sig_x(0), A3 => gl_gr_lg_lh_sig_edges, ZN => gl_gr_lg_lh_n_5);
  gl_gr_lg_lh_g477 : AOI31D0BWP7T port map(A1 => gl_sig_x(2), A2 => gl_sig_x(3), A3 => gl_sig_x(1), B => FE_OFN31_reset, ZN => gl_gr_lg_lh_n_4);
  gl_gr_lg_lh_g478 : NR2D1BWP7T port map(A1 => gl_gr_lg_lh_sig_edges, A2 => FE_OFN31_reset, ZN => gl_gr_lg_lh_n_3);
  gl_gr_lg_lh_count_h_reg_1 : DFD1BWP7T port map(CP => CTS_288, D => gl_gr_lg_lh_n_11, Q => gl_sig_x(1), QN => gl_gr_lg_lh_n_2);
  gl_gr_lg_lh_count_h_reg_0 : DFD1BWP7T port map(CP => CTS_288, D => FE_PHN407_gl_gr_lg_lh_n_9, Q => gl_sig_x(0), QN => gl_gr_lg_lh_n_1);
  gl_gr_lg_lh_count_h_reg_2 : DFD1BWP7T port map(CP => CTS_288, D => FE_PHN406_gl_gr_lg_lh_n_14, Q => gl_sig_x(2), QN => gl_gr_lg_lh_n_0);
  gl_gr_lg_lh_l_edge_g12 : NR2XD0BWP7T port map(A1 => gl_gr_lg_lh_l_edge_n_0, A2 => gl_gr_lg_lh_l_edge_reg2, ZN => gl_gr_lg_lh_sig_edges);
  gl_gr_lg_lh_l_edge_reg2_reg : DFQD1BWP7T port map(CP => CTS_288, D => FE_PHN365_gl_gr_lg_lh_l_edge_reg1, Q => gl_gr_lg_lh_l_edge_reg2);
  gl_gr_lg_lh_l_edge_reg1_reg : DFD1BWP7T port map(CP => CTS_288, D => FE_PHN413_gl_sig_scale_h, Q => gl_gr_lg_lh_l_edge_reg1, QN => gl_gr_lg_lh_l_edge_n_0);
  gl_rom_rom_colour_out_reg_0 : LHQD1BWP7T port map(D => gl_rom_n_1500, E => CTS_322, Q => gl_sig_rom(0));
  gl_rom_rom_colour_out_reg_1 : LHQD1BWP7T port map(D => gl_rom_n_1499, E => CTS_322, Q => gl_sig_rom(1));
  gl_rom_g35179 : MOAI22D0BWP7T port map(A1 => gl_rom_n_1496, A2 => gl_sig_e(9), B1 => gl_rom_n_1498, B2 => gl_sig_e(9), ZN => gl_rom_n_1500);
  gl_rom_g35180 : MOAI22D0BWP7T port map(A1 => gl_rom_n_1497, A2 => gl_sig_e(9), B1 => gl_rom_n_1495, B2 => gl_sig_e(9), ZN => gl_rom_n_1499);
  gl_rom_g35181 : ND4D0BWP7T port map(A1 => gl_rom_n_1490, A2 => gl_rom_n_1488, A3 => gl_rom_n_1481, A4 => gl_rom_n_1480, ZN => gl_rom_n_1498);
  gl_rom_g35182 : AN4D0BWP7T port map(A1 => gl_rom_n_1484, A2 => gl_rom_n_1487, A3 => gl_rom_n_1485, A4 => gl_rom_n_1492, Z => gl_rom_n_1497);
  gl_rom_g35183 : AN4D0BWP7T port map(A1 => gl_rom_n_1493, A2 => gl_rom_n_1494, A3 => gl_rom_n_1486, A4 => gl_rom_n_1482, Z => gl_rom_n_1496);
  gl_rom_g35184 : ND4D0BWP7T port map(A1 => gl_rom_n_1491, A2 => gl_rom_n_1479, A3 => gl_rom_n_1489, A4 => gl_rom_n_1483, ZN => gl_rom_n_1495);
  gl_rom_g35185 : AOI22D0BWP7T port map(A1 => gl_rom_n_1474, A2 => gl_rom_n_38, B1 => gl_rom_n_1463, B2 => gl_rom_n_34, ZN => gl_rom_n_1494);
  gl_rom_g35186 : AOI22D0BWP7T port map(A1 => gl_rom_n_1465, A2 => gl_rom_n_37, B1 => gl_rom_n_1471, B2 => gl_rom_n_31, ZN => gl_rom_n_1493);
  gl_rom_g35187 : AOI22D0BWP7T port map(A1 => gl_rom_n_1469, A2 => gl_rom_n_37, B1 => gl_rom_n_1472, B2 => gl_rom_n_31, ZN => gl_rom_n_1492);
  gl_rom_g35188 : AOI22D0BWP7T port map(A1 => gl_rom_n_1476, A2 => gl_rom_n_37, B1 => gl_rom_n_1462, B2 => gl_rom_n_31, ZN => gl_rom_n_1491);
  gl_rom_g35189 : AOI22D0BWP7T port map(A1 => gl_rom_n_1448, A2 => gl_rom_n_37, B1 => gl_rom_n_1468, B2 => gl_rom_n_31, ZN => gl_rom_n_1490);
  gl_rom_g35190 : AOI22D0BWP7T port map(A1 => gl_rom_n_1473, A2 => gl_rom_n_32, B1 => gl_rom_n_1475, B2 => gl_rom_n_35, ZN => gl_rom_n_1489);
  gl_rom_g35191 : AOI22D0BWP7T port map(A1 => gl_rom_n_1447, A2 => gl_rom_n_32, B1 => gl_rom_n_1470, B2 => gl_rom_n_35, ZN => gl_rom_n_1488);
  gl_rom_g35192 : AOI22D0BWP7T port map(A1 => gl_rom_n_1464, A2 => gl_rom_n_38, B1 => gl_rom_n_1466, B2 => gl_rom_n_34, ZN => gl_rom_n_1487);
  gl_rom_g35193 : AOI22D0BWP7T port map(A1 => gl_rom_n_1450, A2 => gl_rom_n_33, B1 => gl_rom_n_1455, B2 => gl_rom_n_36, ZN => gl_rom_n_1486);
  gl_rom_g35194 : AOI22D0BWP7T port map(A1 => gl_rom_n_1460, A2 => gl_rom_n_33, B1 => gl_rom_n_1478, B2 => gl_rom_n_36, ZN => gl_rom_n_1485);
  gl_rom_g35195 : AOI22D0BWP7T port map(A1 => gl_rom_n_1457, A2 => gl_rom_n_32, B1 => gl_rom_n_1458, B2 => gl_rom_n_35, ZN => gl_rom_n_1484);
  gl_rom_g35196 : AOI22D0BWP7T port map(A1 => gl_rom_n_1453, A2 => gl_rom_n_33, B1 => gl_rom_n_1456, B2 => gl_rom_n_36, ZN => gl_rom_n_1483);
  gl_rom_g35197 : AOI22D0BWP7T port map(A1 => gl_rom_n_1459, A2 => gl_rom_n_32, B1 => gl_rom_n_1461, B2 => gl_rom_n_35, ZN => gl_rom_n_1482);
  gl_rom_g35198 : AOI22D0BWP7T port map(A1 => gl_rom_n_1467, A2 => gl_rom_n_33, B1 => gl_rom_n_1452, B2 => gl_rom_n_36, ZN => gl_rom_n_1481);
  gl_rom_g35199 : AOI22D0BWP7T port map(A1 => gl_rom_n_1477, A2 => gl_rom_n_38, B1 => gl_rom_n_1454, B2 => gl_rom_n_34, ZN => gl_rom_n_1480);
  gl_rom_g35200 : AOI22D0BWP7T port map(A1 => gl_rom_n_1449, A2 => gl_rom_n_38, B1 => gl_rom_n_1451, B2 => gl_rom_n_34, ZN => gl_rom_n_1479);
  gl_rom_g35201 : ND4D0BWP7T port map(A1 => gl_rom_n_1368, A2 => gl_rom_n_1367, A3 => gl_rom_n_1364, A4 => gl_rom_n_1430, ZN => gl_rom_n_1478);
  gl_rom_g35202 : ND4D0BWP7T port map(A1 => gl_rom_n_1404, A2 => gl_rom_n_1414, A3 => gl_rom_n_1400, A4 => gl_rom_n_1392, ZN => gl_rom_n_1477);
  gl_rom_g35203 : ND4D0BWP7T port map(A1 => gl_rom_n_1445, A2 => gl_rom_n_1407, A3 => gl_rom_n_1405, A4 => gl_rom_n_1409, ZN => gl_rom_n_1476);
  gl_rom_g35204 : ND4D0BWP7T port map(A1 => gl_rom_n_1398, A2 => gl_rom_n_1401, A3 => gl_rom_n_1403, A4 => gl_rom_n_1442, ZN => gl_rom_n_1475);
  gl_rom_g35205 : ND4D0BWP7T port map(A1 => gl_rom_n_1443, A2 => gl_rom_n_1399, A3 => gl_rom_n_1395, A4 => gl_rom_n_1391, ZN => gl_rom_n_1474);
  gl_rom_g35206 : ND4D0BWP7T port map(A1 => gl_rom_n_1396, A2 => gl_rom_n_1390, A3 => gl_rom_n_1394, A4 => gl_rom_n_1441, ZN => gl_rom_n_1473);
  gl_rom_g35207 : ND4D0BWP7T port map(A1 => gl_rom_n_1386, A2 => gl_rom_n_1389, A3 => gl_rom_n_1388, A4 => gl_rom_n_1440, ZN => gl_rom_n_1472);
  gl_rom_g35208 : ND4D0BWP7T port map(A1 => gl_rom_n_1387, A2 => gl_rom_n_1439, A3 => gl_rom_n_1381, A4 => gl_rom_n_1385, ZN => gl_rom_n_1471);
  gl_rom_g35209 : ND4D0BWP7T port map(A1 => gl_rom_n_1366, A2 => gl_rom_n_1375, A3 => gl_rom_n_1350, A4 => gl_rom_n_1438, ZN => gl_rom_n_1470);
  gl_rom_g35210 : ND4D0BWP7T port map(A1 => gl_rom_n_1383, A2 => gl_rom_n_1384, A3 => gl_rom_n_1437, A4 => gl_rom_n_1380, ZN => gl_rom_n_1469);
  gl_rom_g35211 : ND4D0BWP7T port map(A1 => gl_rom_n_1422, A2 => gl_rom_n_1349, A3 => gl_rom_n_1402, A4 => gl_rom_n_1363, ZN => gl_rom_n_1468);
  gl_rom_g35212 : ND4D0BWP7T port map(A1 => gl_rom_n_1436, A2 => gl_rom_n_1374, A3 => gl_rom_n_1341, A4 => gl_rom_n_1356, ZN => gl_rom_n_1467);
  gl_rom_g35213 : ND4D0BWP7T port map(A1 => gl_rom_n_1435, A2 => gl_rom_n_1376, A3 => gl_rom_n_1377, A4 => gl_rom_n_1379, ZN => gl_rom_n_1466);
  gl_rom_g35214 : ND4D0BWP7T port map(A1 => gl_rom_n_1378, A2 => gl_rom_n_1434, A3 => gl_rom_n_1369, A4 => gl_rom_n_1372, ZN => gl_rom_n_1465);
  gl_rom_g35215 : ND4D0BWP7T port map(A1 => gl_rom_n_1432, A2 => gl_rom_n_1370, A3 => gl_rom_n_1371, A4 => gl_rom_n_1373, ZN => gl_rom_n_1464);
  gl_rom_g35216 : ND4D0BWP7T port map(A1 => gl_rom_n_1446, A2 => gl_rom_n_1411, A3 => gl_rom_n_1444, A4 => gl_rom_n_1406, ZN => gl_rom_n_1463);
  gl_rom_g35217 : ND4D0BWP7T port map(A1 => gl_rom_n_1412, A2 => gl_rom_n_1410, A3 => gl_rom_n_1413, A4 => gl_rom_n_1415, ZN => gl_rom_n_1462);
  gl_rom_g35218 : ND4D0BWP7T port map(A1 => gl_rom_n_1365, A2 => gl_rom_n_1361, A3 => gl_rom_n_1431, A4 => gl_rom_n_1358, ZN => gl_rom_n_1461);
  gl_rom_g35219 : ND4D0BWP7T port map(A1 => gl_rom_n_1362, A2 => gl_rom_n_1360, A3 => gl_rom_n_1357, A4 => gl_rom_n_1428, ZN => gl_rom_n_1460);
  gl_rom_g35220 : ND4D0BWP7T port map(A1 => gl_rom_n_1347, A2 => gl_rom_n_1351, A3 => gl_rom_n_1426, A4 => gl_rom_n_1344, ZN => gl_rom_n_1459);
  gl_rom_g35221 : ND4D0BWP7T port map(A1 => gl_rom_n_1427, A2 => gl_rom_n_1382, A3 => gl_rom_n_1353, A4 => gl_rom_n_1355, ZN => gl_rom_n_1458);
  gl_rom_g35222 : ND4D0BWP7T port map(A1 => gl_rom_n_1346, A2 => gl_rom_n_1343, A3 => gl_rom_n_1425, A4 => gl_rom_n_1348, ZN => gl_rom_n_1457);
  gl_rom_g35223 : ND4D0BWP7T port map(A1 => gl_rom_n_1342, A2 => gl_rom_n_1340, A3 => gl_rom_n_1423, A4 => gl_rom_n_1338, ZN => gl_rom_n_1456);
  gl_rom_g35224 : ND4D0BWP7T port map(A1 => gl_rom_n_1424, A2 => gl_rom_n_1339, A3 => gl_rom_n_1334, A4 => gl_rom_n_1332, ZN => gl_rom_n_1455);
  gl_rom_g35225 : ND4D0BWP7T port map(A1 => gl_rom_n_1333, A2 => gl_rom_n_1337, A3 => gl_rom_n_1418, A4 => gl_rom_n_1321, ZN => gl_rom_n_1454);
  gl_rom_g35226 : ND4D0BWP7T port map(A1 => gl_rom_n_1335, A2 => gl_rom_n_1331, A3 => gl_rom_n_1421, A4 => gl_rom_n_1336, ZN => gl_rom_n_1453);
  gl_rom_g35227 : ND4D0BWP7T port map(A1 => gl_rom_n_1420, A2 => gl_rom_n_1408, A3 => gl_rom_n_1322, A4 => gl_rom_n_1393, ZN => gl_rom_n_1452);
  gl_rom_g35228 : ND4D0BWP7T port map(A1 => gl_rom_n_1419, A2 => gl_rom_n_1330, A3 => gl_rom_n_1328, A4 => gl_rom_n_1326, ZN => gl_rom_n_1451);
  gl_rom_g35229 : ND4D0BWP7T port map(A1 => gl_rom_n_1327, A2 => gl_rom_n_1329, A3 => gl_rom_n_1320, A4 => gl_rom_n_1416, ZN => gl_rom_n_1450);
  gl_rom_g35230 : ND4D0BWP7T port map(A1 => gl_rom_n_1417, A2 => gl_rom_n_1324, A3 => gl_rom_n_1319, A4 => gl_rom_n_1325, ZN => gl_rom_n_1449);
  gl_rom_g35231 : ND4D0BWP7T port map(A1 => gl_rom_n_1397, A2 => gl_rom_n_1323, A3 => gl_rom_n_1433, A4 => gl_rom_n_1354, ZN => gl_rom_n_1448);
  gl_rom_g35232 : ND4D0BWP7T port map(A1 => gl_rom_n_1345, A2 => gl_rom_n_1359, A3 => gl_rom_n_1352, A4 => gl_rom_n_1429, ZN => gl_rom_n_1447);
  gl_rom_g35233 : AOI22D0BWP7T port map(A1 => gl_rom_n_1312, A2 => gl_rom_n_23, B1 => gl_rom_n_1314, B2 => gl_rom_n_30, ZN => gl_rom_n_1446);
  gl_rom_g35234 : AOI22D0BWP7T port map(A1 => gl_rom_n_1302, A2 => gl_rom_n_25, B1 => gl_rom_n_1303, B2 => gl_rom_n_28, ZN => gl_rom_n_1445);
  gl_rom_g35235 : AOI22D0BWP7T port map(A1 => gl_rom_n_1296, A2 => gl_rom_n_25, B1 => gl_rom_n_1299, B2 => gl_rom_n_28, ZN => gl_rom_n_1444);
  gl_rom_g35236 : AOI22D0BWP7T port map(A1 => gl_rom_n_1281, A2 => gl_rom_n_25, B1 => gl_rom_n_1283, B2 => gl_rom_n_28, ZN => gl_rom_n_1443);
  gl_rom_g35237 : AOI22D0BWP7T port map(A1 => gl_rom_n_1279, A2 => gl_rom_n_25, B1 => gl_rom_n_1280, B2 => gl_rom_n_28, ZN => gl_rom_n_1442);
  gl_rom_g35238 : AOI22D0BWP7T port map(A1 => gl_rom_n_1263, A2 => gl_rom_n_25, B1 => gl_rom_n_1266, B2 => gl_rom_n_28, ZN => gl_rom_n_1441);
  gl_rom_g35239 : AOI22D0BWP7T port map(A1 => gl_rom_n_1254, A2 => gl_rom_n_25, B1 => gl_rom_n_1255, B2 => gl_rom_n_28, ZN => gl_rom_n_1440);
  gl_rom_g35240 : AOI22D0BWP7T port map(A1 => gl_rom_n_1249, A2 => gl_rom_n_25, B1 => gl_rom_n_1251, B2 => gl_rom_n_28, ZN => gl_rom_n_1439);
  gl_rom_g35241 : AOI22D0BWP7T port map(A1 => gl_rom_n_1238, A2 => gl_rom_n_25, B1 => gl_rom_n_1243, B2 => gl_rom_n_28, ZN => gl_rom_n_1438);
  gl_rom_g35242 : AOI22D0BWP7T port map(A1 => gl_rom_n_1239, A2 => gl_rom_n_25, B1 => gl_rom_n_1241, B2 => gl_rom_n_28, ZN => gl_rom_n_1437);
  gl_rom_g35243 : AOI22D0BWP7T port map(A1 => gl_rom_n_1214, A2 => gl_rom_n_25, B1 => gl_rom_n_1223, B2 => gl_rom_n_28, ZN => gl_rom_n_1436);
  gl_rom_g35244 : AOI22D0BWP7T port map(A1 => gl_rom_n_1224, A2 => gl_rom_n_25, B1 => gl_rom_n_1225, B2 => gl_rom_n_28, ZN => gl_rom_n_1435);
  gl_rom_g35245 : AOI22D0BWP7T port map(A1 => gl_rom_n_1218, A2 => gl_rom_n_25, B1 => gl_rom_n_1221, B2 => gl_rom_n_28, ZN => gl_rom_n_1434);
  gl_rom_g35246 : AOI22D0BWP7T port map(A1 => gl_rom_n_1170, A2 => gl_rom_n_25, B1 => gl_rom_n_1199, B2 => gl_rom_n_28, ZN => gl_rom_n_1433);
  gl_rom_g35247 : AOI22D0BWP7T port map(A1 => gl_rom_n_1208, A2 => gl_rom_n_25, B1 => gl_rom_n_1210, B2 => gl_rom_n_28, ZN => gl_rom_n_1432);
  gl_rom_g35248 : AOI22D0BWP7T port map(A1 => gl_rom_n_1185, A2 => gl_rom_n_25, B1 => gl_rom_n_1188, B2 => gl_rom_n_28, ZN => gl_rom_n_1431);
  gl_rom_g35249 : AOI22D0BWP7T port map(A1 => gl_rom_n_1184, A2 => gl_rom_n_25, B1 => gl_rom_n_1186, B2 => gl_rom_n_28, ZN => gl_rom_n_1430);
  gl_rom_g35250 : AOI22D0BWP7T port map(A1 => gl_rom_n_1172, A2 => gl_rom_n_25, B1 => gl_rom_n_1180, B2 => gl_rom_n_28, ZN => gl_rom_n_1429);
  gl_rom_g35251 : AOI22D0BWP7T port map(A1 => gl_rom_n_1167, A2 => gl_rom_n_25, B1 => gl_rom_n_1168, B2 => gl_rom_n_28, ZN => gl_rom_n_1428);
  gl_rom_g35252 : AOI22D0BWP7T port map(A1 => gl_rom_n_1159, A2 => gl_rom_n_25, B1 => gl_rom_n_1160, B2 => gl_rom_n_28, ZN => gl_rom_n_1427);
  gl_rom_g35253 : AOI22D0BWP7T port map(A1 => gl_rom_n_1153, A2 => gl_rom_n_25, B1 => gl_rom_n_1157, B2 => gl_rom_n_28, ZN => gl_rom_n_1426);
  gl_rom_g35254 : AOI22D0BWP7T port map(A1 => gl_rom_n_1144, A2 => gl_rom_n_25, B1 => gl_rom_n_1145, B2 => gl_rom_n_28, ZN => gl_rom_n_1425);
  gl_rom_g35255 : AOI22D0BWP7T port map(A1 => gl_rom_n_1121, A2 => gl_rom_n_25, B1 => gl_rom_n_1123, B2 => gl_rom_n_28, ZN => gl_rom_n_1424);
  gl_rom_g35256 : AOI22D0BWP7T port map(A1 => gl_rom_n_1119, A2 => gl_rom_n_25, B1 => gl_rom_n_1120, B2 => gl_rom_n_28, ZN => gl_rom_n_1423);
  gl_rom_g35257 : AOI22D0BWP7T port map(A1 => gl_rom_n_1191, A2 => gl_rom_n_25, B1 => gl_rom_n_1084, B2 => gl_rom_n_28, ZN => gl_rom_n_1422);
  gl_rom_g35258 : AOI22D0BWP7T port map(A1 => gl_rom_n_1103, A2 => gl_rom_n_25, B1 => gl_rom_n_1104, B2 => gl_rom_n_28, ZN => gl_rom_n_1421);
  gl_rom_g35259 : AOI22D0BWP7T port map(A1 => gl_rom_n_1085, A2 => gl_rom_n_25, B1 => gl_rom_n_1101, B2 => gl_rom_n_28, ZN => gl_rom_n_1420);
  gl_rom_g35260 : AOI22D0BWP7T port map(A1 => gl_rom_n_1095, A2 => gl_rom_n_25, B1 => gl_rom_n_1097, B2 => gl_rom_n_28, ZN => gl_rom_n_1419);
  gl_rom_g35261 : AOI22D0BWP7T port map(A1 => gl_rom_n_1076, A2 => gl_rom_n_25, B1 => gl_rom_n_1082, B2 => gl_rom_n_28, ZN => gl_rom_n_1418);
  gl_rom_g35262 : AOI22D0BWP7T port map(A1 => gl_rom_n_1078, A2 => gl_rom_n_25, B1 => gl_rom_n_1079, B2 => gl_rom_n_28, ZN => gl_rom_n_1417);
  gl_rom_g35263 : AOI22D0BWP7T port map(A1 => gl_rom_n_1073, A2 => gl_rom_n_25, B1 => gl_rom_n_1075, B2 => gl_rom_n_28, ZN => gl_rom_n_1416);
  gl_rom_g35264 : AOI22D0BWP7T port map(A1 => gl_rom_n_1317, A2 => gl_rom_n_25, B1 => gl_rom_n_1190, B2 => gl_rom_n_28, ZN => gl_rom_n_1415);
  gl_rom_g35265 : AOI22D0BWP7T port map(A1 => gl_rom_n_1300, A2 => gl_rom_n_25, B1 => gl_rom_n_1306, B2 => gl_rom_n_28, ZN => gl_rom_n_1414);
  gl_rom_g35266 : AOI22D0BWP7T port map(A1 => gl_rom_n_1313, A2 => gl_rom_n_26, B1 => gl_rom_n_1316, B2 => gl_rom_n_27, ZN => gl_rom_n_1413);
  gl_rom_g35267 : AOI22D0BWP7T port map(A1 => gl_rom_n_1309, A2 => gl_rom_n_23, B1 => gl_rom_n_1311, B2 => gl_rom_n_30, ZN => gl_rom_n_1412);
  gl_rom_g35268 : AOI22D0BWP7T port map(A1 => gl_rom_n_1304, A2 => gl_rom_n_26, B1 => gl_rom_n_1307, B2 => gl_rom_n_27, ZN => gl_rom_n_1411);
  gl_rom_g35269 : AOI22D0BWP7T port map(A1 => gl_rom_n_1305, A2 => gl_rom_n_24, B1 => gl_rom_n_1308, B2 => gl_rom_n_29, ZN => gl_rom_n_1410);
  gl_rom_g35270 : AOI22D0BWP7T port map(A1 => gl_rom_n_1298, A2 => gl_rom_n_23, B1 => gl_rom_n_1301, B2 => gl_rom_n_30, ZN => gl_rom_n_1409);
  gl_rom_g35271 : AOI22D0BWP7T port map(A1 => gl_rom_n_1277, A2 => gl_rom_n_26, B1 => gl_rom_n_1294, B2 => gl_rom_n_27, ZN => gl_rom_n_1408);
  gl_rom_g35272 : AOI22D0BWP7T port map(A1 => gl_rom_n_1295, A2 => gl_rom_n_26, B1 => gl_rom_n_1297, B2 => gl_rom_n_27, ZN => gl_rom_n_1407);
  gl_rom_g35273 : AOI22D0BWP7T port map(A1 => gl_rom_n_1288, A2 => gl_rom_n_24, B1 => gl_rom_n_1291, B2 => gl_rom_n_29, ZN => gl_rom_n_1406);
  gl_rom_g35274 : AOI22D0BWP7T port map(A1 => gl_rom_n_1289, A2 => gl_rom_n_24, B1 => gl_rom_n_1293, B2 => gl_rom_n_29, ZN => gl_rom_n_1405);
  gl_rom_g35275 : AOI22D0BWP7T port map(A1 => gl_rom_n_1284, A2 => gl_rom_n_23, B1 => gl_rom_n_1290, B2 => gl_rom_n_30, ZN => gl_rom_n_1404);
  gl_rom_g35276 : AOI22D0BWP7T port map(A1 => gl_rom_n_1286, A2 => gl_rom_n_23, B1 => gl_rom_n_1287, B2 => gl_rom_n_30, ZN => gl_rom_n_1403);
  gl_rom_g35277 : AOI22D0BWP7T port map(A1 => gl_rom_n_1200, A2 => gl_rom_n_26, B1 => gl_rom_n_1264, B2 => gl_rom_n_27, ZN => gl_rom_n_1402);
  gl_rom_g35278 : AOI22D0BWP7T port map(A1 => gl_rom_n_1282, A2 => gl_rom_n_26, B1 => gl_rom_n_1285, B2 => gl_rom_n_27, ZN => gl_rom_n_1401);
  gl_rom_g35279 : AOI22D0BWP7T port map(A1 => gl_rom_n_1267, A2 => gl_rom_n_26, B1 => gl_rom_n_1275, B2 => gl_rom_n_27, ZN => gl_rom_n_1400);
  gl_rom_g35280 : AOI22D0BWP7T port map(A1 => gl_rom_n_1273, A2 => gl_rom_n_26, B1 => gl_rom_n_1276, B2 => gl_rom_n_27, ZN => gl_rom_n_1399);
  gl_rom_g35281 : AOI22D0BWP7T port map(A1 => gl_rom_n_1274, A2 => gl_rom_n_24, B1 => gl_rom_n_1278, B2 => gl_rom_n_29, ZN => gl_rom_n_1398);
  gl_rom_g35282 : AOI22D0BWP7T port map(A1 => gl_rom_n_1231, A2 => gl_rom_n_26, B1 => gl_rom_n_1262, B2 => gl_rom_n_27, ZN => gl_rom_n_1397);
  gl_rom_g35283 : AOI22D0BWP7T port map(A1 => gl_rom_n_1271, A2 => gl_rom_n_23, B1 => gl_rom_n_1272, B2 => gl_rom_n_30, ZN => gl_rom_n_1396);
  gl_rom_g35284 : AOI22D0BWP7T port map(A1 => gl_rom_n_1265, A2 => gl_rom_n_23, B1 => gl_rom_n_1269, B2 => gl_rom_n_30, ZN => gl_rom_n_1395);
  gl_rom_g35285 : AOI22D0BWP7T port map(A1 => gl_rom_n_1268, A2 => gl_rom_n_26, B1 => gl_rom_n_1270, B2 => gl_rom_n_27, ZN => gl_rom_n_1394);
  gl_rom_g35286 : AOI22D0BWP7T port map(A1 => gl_rom_n_1245, A2 => gl_rom_n_24, B1 => gl_rom_n_1261, B2 => gl_rom_n_29, ZN => gl_rom_n_1393);
  gl_rom_g35287 : AOI22D0BWP7T port map(A1 => gl_rom_n_1253, A2 => gl_rom_n_24, B1 => gl_rom_n_1259, B2 => gl_rom_n_29, ZN => gl_rom_n_1392);
  gl_rom_g35288 : AOI22D0BWP7T port map(A1 => gl_rom_n_1256, A2 => gl_rom_n_24, B1 => gl_rom_n_1258, B2 => gl_rom_n_29, ZN => gl_rom_n_1391);
  gl_rom_g35289 : AOI22D0BWP7T port map(A1 => gl_rom_n_1257, A2 => gl_rom_n_24, B1 => gl_rom_n_1260, B2 => gl_rom_n_29, ZN => gl_rom_n_1390);
  gl_rom_g35290 : AOI22D0BWP7T port map(A1 => gl_rom_n_1250, A2 => gl_rom_n_26, B1 => gl_rom_n_1252, B2 => gl_rom_n_27, ZN => gl_rom_n_1389);
  gl_rom_g35291 : AOI22D0BWP7T port map(A1 => gl_rom_n_1247, A2 => gl_rom_n_23, B1 => gl_rom_n_1248, B2 => gl_rom_n_30, ZN => gl_rom_n_1388);
  gl_rom_g35292 : AOI22D0BWP7T port map(A1 => gl_rom_n_1240, A2 => gl_rom_n_26, B1 => gl_rom_n_1244, B2 => gl_rom_n_27, ZN => gl_rom_n_1387);
  gl_rom_g35293 : AOI22D0BWP7T port map(A1 => gl_rom_n_1242, A2 => gl_rom_n_24, B1 => gl_rom_n_1246, B2 => gl_rom_n_29, ZN => gl_rom_n_1386);
  gl_rom_g35294 : AOI22D0BWP7T port map(A1 => gl_rom_n_1234, A2 => gl_rom_n_23, B1 => gl_rom_n_1236, B2 => gl_rom_n_30, ZN => gl_rom_n_1385);
  gl_rom_g35295 : AOI22D0BWP7T port map(A1 => gl_rom_n_1235, A2 => gl_rom_n_26, B1 => gl_rom_n_1237, B2 => gl_rom_n_27, ZN => gl_rom_n_1384);
  gl_rom_g35296 : AOI22D0BWP7T port map(A1 => gl_rom_n_1232, A2 => gl_rom_n_23, B1 => gl_rom_n_1233, B2 => gl_rom_n_30, ZN => gl_rom_n_1383);
  gl_rom_g35297 : AOI22D0BWP7T port map(A1 => gl_rom_n_1147, A2 => gl_rom_n_24, B1 => gl_rom_n_1150, B2 => gl_rom_n_29, ZN => gl_rom_n_1382);
  gl_rom_g35298 : AOI22D0BWP7T port map(A1 => gl_rom_n_1226, A2 => gl_rom_n_24, B1 => gl_rom_n_1229, B2 => gl_rom_n_29, ZN => gl_rom_n_1381);
  gl_rom_g35299 : AOI22D0BWP7T port map(A1 => gl_rom_n_1228, A2 => gl_rom_n_24, B1 => gl_rom_n_1230, B2 => gl_rom_n_29, ZN => gl_rom_n_1380);
  gl_rom_g35300 : AOI22D0BWP7T port map(A1 => gl_rom_n_1219, A2 => gl_rom_n_23, B1 => gl_rom_n_1222, B2 => gl_rom_n_30, ZN => gl_rom_n_1379);
  gl_rom_g35301 : AOI22D0BWP7T port map(A1 => gl_rom_n_1209, A2 => gl_rom_n_23, B1 => gl_rom_n_1213, B2 => gl_rom_n_30, ZN => gl_rom_n_1378);
  gl_rom_g35302 : AOI22D0BWP7T port map(A1 => gl_rom_n_1216, A2 => gl_rom_n_26, B1 => gl_rom_n_1217, B2 => gl_rom_n_27, ZN => gl_rom_n_1377);
  gl_rom_g35303 : AOI22D0BWP7T port map(A1 => gl_rom_n_1211, A2 => gl_rom_n_24, B1 => gl_rom_n_1215, B2 => gl_rom_n_29, ZN => gl_rom_n_1376);
  gl_rom_g35304 : AOI22D0BWP7T port map(A1 => gl_rom_n_1207, A2 => gl_rom_n_26, B1 => gl_rom_n_1212, B2 => gl_rom_n_27, ZN => gl_rom_n_1375);
  gl_rom_g35305 : AOI22D0BWP7T port map(A1 => gl_rom_n_1183, A2 => gl_rom_n_23, B1 => gl_rom_n_1197, B2 => gl_rom_n_30, ZN => gl_rom_n_1374);
  gl_rom_g35306 : AOI22D0BWP7T port map(A1 => gl_rom_n_1204, A2 => gl_rom_n_23, B1 => gl_rom_n_1206, B2 => gl_rom_n_30, ZN => gl_rom_n_1373);
  gl_rom_g35307 : AOI22D0BWP7T port map(A1 => gl_rom_n_1203, A2 => gl_rom_n_26, B1 => gl_rom_n_1205, B2 => gl_rom_n_27, ZN => gl_rom_n_1372);
  gl_rom_g35308 : AOI22D0BWP7T port map(A1 => gl_rom_n_1201, A2 => gl_rom_n_26, B1 => gl_rom_n_1202, B2 => gl_rom_n_27, ZN => gl_rom_n_1371);
  gl_rom_g35309 : AOI22D0BWP7T port map(A1 => gl_rom_n_1194, A2 => gl_rom_n_24, B1 => gl_rom_n_1198, B2 => gl_rom_n_29, ZN => gl_rom_n_1370);
  gl_rom_g35310 : AOI22D0BWP7T port map(A1 => gl_rom_n_1193, A2 => gl_rom_n_24, B1 => gl_rom_n_1196, B2 => gl_rom_n_29, ZN => gl_rom_n_1369);
  gl_rom_g35311 : AOI22D0BWP7T port map(A1 => gl_rom_n_1318, A2 => gl_rom_n_26, B1 => gl_rom_n_1192, B2 => gl_rom_n_27, ZN => gl_rom_n_1368);
  gl_rom_g35312 : AOI22D0BWP7T port map(A1 => gl_rom_n_1187, A2 => gl_rom_n_23, B1 => gl_rom_n_1189, B2 => gl_rom_n_30, ZN => gl_rom_n_1367);
  gl_rom_g35313 : AOI22D0BWP7T port map(A1 => gl_rom_n_1063, A2 => gl_rom_n_24, B1 => gl_rom_n_1195, B2 => gl_rom_n_29, ZN => gl_rom_n_1366);
  gl_rom_g35314 : AOI22D0BWP7T port map(A1 => gl_rom_n_1177, A2 => gl_rom_n_23, B1 => gl_rom_n_1181, B2 => gl_rom_n_30, ZN => gl_rom_n_1365);
  gl_rom_g35315 : AOI22D0BWP7T port map(A1 => gl_rom_n_1179, A2 => gl_rom_n_24, B1 => gl_rom_n_1182, B2 => gl_rom_n_29, ZN => gl_rom_n_1364);
  gl_rom_g35316 : AOI22D0BWP7T port map(A1 => gl_rom_n_1086, A2 => gl_rom_n_23, B1 => gl_rom_n_1178, B2 => gl_rom_n_30, ZN => gl_rom_n_1363);
  gl_rom_g35317 : AOI22D0BWP7T port map(A1 => gl_rom_n_1175, A2 => gl_rom_n_23, B1 => gl_rom_n_1176, B2 => gl_rom_n_30, ZN => gl_rom_n_1362);
  gl_rom_g35318 : AOI22D0BWP7T port map(A1 => gl_rom_n_1169, A2 => gl_rom_n_26, B1 => gl_rom_n_1173, B2 => gl_rom_n_27, ZN => gl_rom_n_1361);
  gl_rom_g35319 : AOI22D0BWP7T port map(A1 => gl_rom_n_1171, A2 => gl_rom_n_26, B1 => gl_rom_n_1174, B2 => gl_rom_n_27, ZN => gl_rom_n_1360);
  gl_rom_g35320 : AOI22D0BWP7T port map(A1 => gl_rom_n_1156, A2 => gl_rom_n_23, B1 => gl_rom_n_1163, B2 => gl_rom_n_30, ZN => gl_rom_n_1359);
  gl_rom_g35321 : AOI22D0BWP7T port map(A1 => gl_rom_n_1161, A2 => gl_rom_n_24, B1 => gl_rom_n_1164, B2 => gl_rom_n_29, ZN => gl_rom_n_1358);
  gl_rom_g35322 : AOI22D0BWP7T port map(A1 => gl_rom_n_1162, A2 => gl_rom_n_24, B1 => gl_rom_n_1166, B2 => gl_rom_n_29, ZN => gl_rom_n_1357);
  gl_rom_g35323 : AOI22D0BWP7T port map(A1 => gl_rom_n_1151, A2 => gl_rom_n_26, B1 => gl_rom_n_1165, B2 => gl_rom_n_27, ZN => gl_rom_n_1356);
  gl_rom_g35324 : AOI22D0BWP7T port map(A1 => gl_rom_n_1155, A2 => gl_rom_n_23, B1 => gl_rom_n_1158, B2 => gl_rom_n_30, ZN => gl_rom_n_1355);
  gl_rom_g35325 : AOI22D0BWP7T port map(A1 => gl_rom_n_1118, A2 => gl_rom_n_24, B1 => gl_rom_n_1135, B2 => gl_rom_n_29, ZN => gl_rom_n_1354);
  gl_rom_g35326 : AOI22D0BWP7T port map(A1 => gl_rom_n_1152, A2 => gl_rom_n_26, B1 => gl_rom_n_1154, B2 => gl_rom_n_27, ZN => gl_rom_n_1353);
  gl_rom_g35327 : AOI22D0BWP7T port map(A1 => gl_rom_n_1143, A2 => gl_rom_n_26, B1 => gl_rom_n_1148, B2 => gl_rom_n_27, ZN => gl_rom_n_1352);
  gl_rom_g35328 : AOI22D0BWP7T port map(A1 => gl_rom_n_1146, A2 => gl_rom_n_23, B1 => gl_rom_n_1149, B2 => gl_rom_n_30, ZN => gl_rom_n_1351);
  gl_rom_g35329 : AOI22D0BWP7T port map(A1 => gl_rom_n_1220, A2 => gl_rom_n_23, B1 => gl_rom_n_1227, B2 => gl_rom_n_30, ZN => gl_rom_n_1350);
  gl_rom_g35330 : AOI22D0BWP7T port map(A1 => gl_rom_n_1109, A2 => gl_rom_n_24, B1 => gl_rom_n_1139, B2 => gl_rom_n_29, ZN => gl_rom_n_1349);
  gl_rom_g35331 : AOI22D0BWP7T port map(A1 => gl_rom_n_1140, A2 => gl_rom_n_26, B1 => gl_rom_n_1142, B2 => gl_rom_n_27, ZN => gl_rom_n_1348);
  gl_rom_g35332 : AOI22D0BWP7T port map(A1 => gl_rom_n_1138, A2 => gl_rom_n_26, B1 => gl_rom_n_1141, B2 => gl_rom_n_27, ZN => gl_rom_n_1347);
  gl_rom_g35333 : AOI22D0BWP7T port map(A1 => gl_rom_n_1136, A2 => gl_rom_n_23, B1 => gl_rom_n_1137, B2 => gl_rom_n_30, ZN => gl_rom_n_1346);
  gl_rom_g35334 : AOI22D0BWP7T port map(A1 => gl_rom_n_1128, A2 => gl_rom_n_24, B1 => gl_rom_n_1131, B2 => gl_rom_n_29, ZN => gl_rom_n_1345);
  gl_rom_g35335 : AOI22D0BWP7T port map(A1 => gl_rom_n_1129, A2 => gl_rom_n_24, B1 => gl_rom_n_1132, B2 => gl_rom_n_29, ZN => gl_rom_n_1344);
  gl_rom_g35336 : AOI22D0BWP7T port map(A1 => gl_rom_n_1130, A2 => gl_rom_n_24, B1 => gl_rom_n_1134, B2 => gl_rom_n_29, ZN => gl_rom_n_1343);
  gl_rom_g35337 : AOI22D0BWP7T port map(A1 => gl_rom_n_1126, A2 => gl_rom_n_23, B1 => gl_rom_n_1127, B2 => gl_rom_n_30, ZN => gl_rom_n_1342);
  gl_rom_g35338 : AOI22D0BWP7T port map(A1 => gl_rom_n_1125, A2 => gl_rom_n_24, B1 => gl_rom_n_1133, B2 => gl_rom_n_29, ZN => gl_rom_n_1341);
  gl_rom_g35339 : AOI22D0BWP7T port map(A1 => gl_rom_n_1122, A2 => gl_rom_n_26, B1 => gl_rom_n_1124, B2 => gl_rom_n_27, ZN => gl_rom_n_1340);
  gl_rom_g35340 : AOI22D0BWP7T port map(A1 => gl_rom_n_1113, A2 => gl_rom_n_23, B1 => gl_rom_n_1116, B2 => gl_rom_n_30, ZN => gl_rom_n_1339);
  gl_rom_g35341 : AOI22D0BWP7T port map(A1 => gl_rom_n_1114, A2 => gl_rom_n_24, B1 => gl_rom_n_1117, B2 => gl_rom_n_29, ZN => gl_rom_n_1338);
  gl_rom_g35342 : AOI22D0BWP7T port map(A1 => gl_rom_n_1107, A2 => gl_rom_n_23, B1 => gl_rom_n_1115, B2 => gl_rom_n_30, ZN => gl_rom_n_1337);
  gl_rom_g35343 : AOI22D0BWP7T port map(A1 => gl_rom_n_1111, A2 => gl_rom_n_26, B1 => gl_rom_n_1112, B2 => gl_rom_n_27, ZN => gl_rom_n_1336);
  gl_rom_g35344 : AOI22D0BWP7T port map(A1 => gl_rom_n_1106, A2 => gl_rom_n_23, B1 => gl_rom_n_1110, B2 => gl_rom_n_30, ZN => gl_rom_n_1335);
  gl_rom_g35345 : AOI22D0BWP7T port map(A1 => gl_rom_n_1105, A2 => gl_rom_n_26, B1 => gl_rom_n_1108, B2 => gl_rom_n_27, ZN => gl_rom_n_1334);
  gl_rom_g35346 : AOI22D0BWP7T port map(A1 => gl_rom_n_1094, A2 => gl_rom_n_26, B1 => gl_rom_n_1099, B2 => gl_rom_n_27, ZN => gl_rom_n_1333);
  gl_rom_g35347 : AOI22D0BWP7T port map(A1 => gl_rom_n_1096, A2 => gl_rom_n_24, B1 => gl_rom_n_1100, B2 => gl_rom_n_29, ZN => gl_rom_n_1332);
  gl_rom_g35348 : AOI22D0BWP7T port map(A1 => gl_rom_n_1098, A2 => gl_rom_n_24, B1 => gl_rom_n_1102, B2 => gl_rom_n_29, ZN => gl_rom_n_1331);
  gl_rom_g35349 : AOI22D0BWP7T port map(A1 => gl_rom_n_1091, A2 => gl_rom_n_26, B1 => gl_rom_n_1093, B2 => gl_rom_n_27, ZN => gl_rom_n_1330);
  gl_rom_g35350 : AOI22D0BWP7T port map(A1 => gl_rom_n_1090, A2 => gl_rom_n_26, B1 => gl_rom_n_1092, B2 => gl_rom_n_27, ZN => gl_rom_n_1329);
  gl_rom_g35351 : AOI22D0BWP7T port map(A1 => gl_rom_n_1088, A2 => gl_rom_n_23, B1 => gl_rom_n_1089, B2 => gl_rom_n_30, ZN => gl_rom_n_1328);
  gl_rom_g35352 : AOI22D0BWP7T port map(A1 => gl_rom_n_1080, A2 => gl_rom_n_23, B1 => gl_rom_n_1083, B2 => gl_rom_n_30, ZN => gl_rom_n_1327);
  gl_rom_g35353 : AOI22D0BWP7T port map(A1 => gl_rom_n_1081, A2 => gl_rom_n_24, B1 => gl_rom_n_1087, B2 => gl_rom_n_29, ZN => gl_rom_n_1326);
  gl_rom_g35354 : AOI22D0BWP7T port map(A1 => gl_rom_n_1074, A2 => gl_rom_n_26, B1 => gl_rom_n_1077, B2 => gl_rom_n_27, ZN => gl_rom_n_1325);
  gl_rom_g35355 : AOI22D0BWP7T port map(A1 => gl_rom_n_1071, A2 => gl_rom_n_23, B1 => gl_rom_n_1072, B2 => gl_rom_n_30, ZN => gl_rom_n_1324);
  gl_rom_g35356 : AOI22D0BWP7T port map(A1 => gl_rom_n_1292, A2 => gl_rom_n_23, B1 => gl_rom_n_1065, B2 => gl_rom_n_30, ZN => gl_rom_n_1323);
  gl_rom_g35357 : AOI22D0BWP7T port map(A1 => gl_rom_n_1310, A2 => gl_rom_n_23, B1 => gl_rom_n_1070, B2 => gl_rom_n_30, ZN => gl_rom_n_1322);
  gl_rom_g35358 : AOI22D0BWP7T port map(A1 => gl_rom_n_1315, A2 => gl_rom_n_24, B1 => gl_rom_n_1067, B2 => gl_rom_n_29, ZN => gl_rom_n_1321);
  gl_rom_g35359 : AOI22D0BWP7T port map(A1 => gl_rom_n_1064, A2 => gl_rom_n_24, B1 => gl_rom_n_1068, B2 => gl_rom_n_29, ZN => gl_rom_n_1320);
  gl_rom_g35360 : AOI22D0BWP7T port map(A1 => gl_rom_n_1066, A2 => gl_rom_n_24, B1 => gl_rom_n_1069, B2 => gl_rom_n_29, ZN => gl_rom_n_1319);
  gl_rom_g35361 : ND4D0BWP7T port map(A1 => gl_rom_n_294, A2 => gl_rom_n_549, A3 => gl_rom_n_546, A4 => gl_rom_n_547, ZN => gl_rom_n_1318);
  gl_rom_g35362 : ND4D0BWP7T port map(A1 => gl_rom_n_1056, A2 => gl_rom_n_1059, A3 => gl_rom_n_1058, A4 => gl_rom_n_1054, ZN => gl_rom_n_1317);
  gl_rom_g35363 : ND4D0BWP7T port map(A1 => gl_rom_n_1052, A2 => gl_rom_n_1048, A3 => gl_rom_n_1047, A4 => gl_rom_n_1051, ZN => gl_rom_n_1316);
  gl_rom_g35364 : ND4D0BWP7T port map(A1 => gl_rom_n_1046, A2 => gl_rom_n_1050, A3 => gl_rom_n_1038, A4 => gl_rom_n_1033, ZN => gl_rom_n_1315);
  gl_rom_g35365 : ND4D0BWP7T port map(A1 => gl_rom_n_1045, A2 => gl_rom_n_1049, A3 => gl_rom_n_1042, A4 => gl_rom_n_1040, ZN => gl_rom_n_1314);
  gl_rom_g35366 : ND4D0BWP7T port map(A1 => gl_rom_n_1039, A2 => gl_rom_n_1044, A3 => gl_rom_n_1041, A4 => gl_rom_n_1043, ZN => gl_rom_n_1313);
  gl_rom_g35367 : ND4D0BWP7T port map(A1 => gl_rom_n_1030, A2 => gl_rom_n_1034, A3 => gl_rom_n_1027, A4 => gl_rom_n_1024, ZN => gl_rom_n_1312);
  gl_rom_g35368 : ND4D0BWP7T port map(A1 => gl_rom_n_1031, A2 => gl_rom_n_1037, A3 => gl_rom_n_1032, A4 => gl_rom_n_1035, ZN => gl_rom_n_1311);
  gl_rom_g35369 : ND4D0BWP7T port map(A1 => gl_rom_n_1010, A2 => gl_rom_n_1020, A3 => gl_rom_n_988, A4 => gl_rom_n_982, ZN => gl_rom_n_1310);
  gl_rom_g35370 : ND4D0BWP7T port map(A1 => gl_rom_n_1023, A2 => gl_rom_n_1029, A3 => gl_rom_n_1025, A4 => gl_rom_n_1028, ZN => gl_rom_n_1309);
  gl_rom_g35371 : ND4D0BWP7T port map(A1 => gl_rom_n_1021, A2 => gl_rom_n_1017, A3 => gl_rom_n_1016, A4 => gl_rom_n_1019, ZN => gl_rom_n_1308);
  gl_rom_g35372 : ND4D0BWP7T port map(A1 => gl_rom_n_1015, A2 => gl_rom_n_1018, A3 => gl_rom_n_1012, A4 => gl_rom_n_1007, ZN => gl_rom_n_1307);
  gl_rom_g35373 : ND4D0BWP7T port map(A1 => gl_rom_n_1005, A2 => gl_rom_n_1014, A3 => gl_rom_n_1000, A4 => gl_rom_n_997, ZN => gl_rom_n_1306);
  gl_rom_g35374 : ND4D0BWP7T port map(A1 => gl_rom_n_1008, A2 => gl_rom_n_1013, A3 => gl_rom_n_1009, A4 => gl_rom_n_1011, ZN => gl_rom_n_1305);
  gl_rom_g35375 : ND4D0BWP7T port map(A1 => gl_rom_n_999, A2 => gl_rom_n_1002, A3 => gl_rom_n_995, A4 => gl_rom_n_990, ZN => gl_rom_n_1304);
  gl_rom_g35376 : ND4D0BWP7T port map(A1 => gl_rom_n_1006, A2 => gl_rom_n_1003, A3 => gl_rom_n_998, A4 => gl_rom_n_1001, ZN => gl_rom_n_1303);
  gl_rom_g35377 : ND4D0BWP7T port map(A1 => gl_rom_n_996, A2 => gl_rom_n_993, A3 => gl_rom_n_994, A4 => gl_rom_n_992, ZN => gl_rom_n_1302);
  gl_rom_g35378 : ND4D0BWP7T port map(A1 => gl_rom_n_986, A2 => gl_rom_n_991, A3 => gl_rom_n_989, A4 => gl_rom_n_984, ZN => gl_rom_n_1301);
  gl_rom_g35379 : ND4D0BWP7T port map(A1 => gl_rom_n_975, A2 => gl_rom_n_985, A3 => gl_rom_n_971, A4 => gl_rom_n_965, ZN => gl_rom_n_1300);
  gl_rom_g35380 : ND4D0BWP7T port map(A1 => gl_rom_n_983, A2 => gl_rom_n_987, A3 => gl_rom_n_979, A4 => gl_rom_n_977, ZN => gl_rom_n_1299);
  gl_rom_g35381 : ND4D0BWP7T port map(A1 => gl_rom_n_978, A2 => gl_rom_n_981, A3 => gl_rom_n_980, A4 => gl_rom_n_976, ZN => gl_rom_n_1298);
  gl_rom_g35382 : ND4D0BWP7T port map(A1 => gl_rom_n_968, A2 => gl_rom_n_974, A3 => gl_rom_n_970, A4 => gl_rom_n_973, ZN => gl_rom_n_1297);
  gl_rom_g35383 : ND4D0BWP7T port map(A1 => gl_rom_n_969, A2 => gl_rom_n_972, A3 => gl_rom_n_964, A4 => gl_rom_n_962, ZN => gl_rom_n_1296);
  gl_rom_g35384 : ND4D0BWP7T port map(A1 => gl_rom_n_967, A2 => gl_rom_n_961, A3 => gl_rom_n_960, A4 => gl_rom_n_963, ZN => gl_rom_n_1295);
  gl_rom_g35385 : ND4D0BWP7T port map(A1 => gl_rom_n_956, A2 => gl_rom_n_928, A3 => gl_rom_n_918, A4 => gl_rom_n_943, ZN => gl_rom_n_1294);
  gl_rom_g35386 : ND4D0BWP7T port map(A1 => gl_rom_n_959, A2 => gl_rom_n_955, A3 => gl_rom_n_958, A4 => gl_rom_n_954, ZN => gl_rom_n_1293);
  gl_rom_g35387 : ND4D0BWP7T port map(A1 => gl_rom_n_899, A2 => gl_rom_n_952, A3 => gl_rom_n_925, A4 => gl_rom_n_867, ZN => gl_rom_n_1292);
  gl_rom_g35388 : ND4D0BWP7T port map(A1 => gl_rom_n_953, A2 => gl_rom_n_957, A3 => gl_rom_n_949, A4 => gl_rom_n_946, ZN => gl_rom_n_1291);
  gl_rom_g35389 : ND4D0BWP7T port map(A1 => gl_rom_n_947, A2 => gl_rom_n_950, A3 => gl_rom_n_939, A4 => gl_rom_n_933, ZN => gl_rom_n_1290);
  gl_rom_g35390 : ND4D0BWP7T port map(A1 => gl_rom_n_945, A2 => gl_rom_n_951, A3 => gl_rom_n_948, A4 => gl_rom_n_944, ZN => gl_rom_n_1289);
  gl_rom_g35391 : ND4D0BWP7T port map(A1 => gl_rom_n_936, A2 => gl_rom_n_941, A3 => gl_rom_n_935, A4 => gl_rom_n_931, ZN => gl_rom_n_1288);
  gl_rom_g35392 : ND4D0BWP7T port map(A1 => gl_rom_n_940, A2 => gl_rom_n_942, A3 => gl_rom_n_938, A4 => gl_rom_n_937, ZN => gl_rom_n_1287);
  gl_rom_g35393 : ND4D0BWP7T port map(A1 => gl_rom_n_932, A2 => gl_rom_n_934, A3 => gl_rom_n_930, A4 => gl_rom_n_929, ZN => gl_rom_n_1286);
  gl_rom_g35394 : ND4D0BWP7T port map(A1 => gl_rom_n_927, A2 => gl_rom_n_926, A3 => gl_rom_n_922, A4 => gl_rom_n_923, ZN => gl_rom_n_1285);
  gl_rom_g35395 : ND4D0BWP7T port map(A1 => gl_rom_n_921, A2 => gl_rom_n_909, A3 => gl_rom_n_902, A4 => gl_rom_n_916, ZN => gl_rom_n_1284);
  gl_rom_g35396 : ND4D0BWP7T port map(A1 => gl_rom_n_914, A2 => gl_rom_n_924, A3 => gl_rom_n_915, A4 => gl_rom_n_920, ZN => gl_rom_n_1283);
  gl_rom_g35397 : ND4D0BWP7T port map(A1 => gl_rom_n_913, A2 => gl_rom_n_919, A3 => gl_rom_n_917, A4 => gl_rom_n_912, ZN => gl_rom_n_1282);
  gl_rom_g35398 : ND4D0BWP7T port map(A1 => gl_rom_n_906, A2 => gl_rom_n_907, A3 => gl_rom_n_901, A4 => gl_rom_n_897, ZN => gl_rom_n_1281);
  gl_rom_g35399 : ND4D0BWP7T port map(A1 => gl_rom_n_911, A2 => gl_rom_n_905, A3 => gl_rom_n_904, A4 => gl_rom_n_908, ZN => gl_rom_n_1280);
  gl_rom_g35400 : ND4D0BWP7T port map(A1 => gl_rom_n_903, A2 => gl_rom_n_898, A3 => gl_rom_n_896, A4 => gl_rom_n_900, ZN => gl_rom_n_1279);
  gl_rom_g35401 : ND4D0BWP7T port map(A1 => gl_rom_n_893, A2 => gl_rom_n_894, A3 => gl_rom_n_891, A4 => gl_rom_n_889, ZN => gl_rom_n_1278);
  gl_rom_g35402 : ND4D0BWP7T port map(A1 => gl_rom_n_895, A2 => gl_rom_n_879, A3 => gl_rom_n_860, A4 => gl_rom_n_863, ZN => gl_rom_n_1277);
  gl_rom_g35403 : ND4D0BWP7T port map(A1 => gl_rom_n_892, A2 => gl_rom_n_885, A3 => gl_rom_n_880, A4 => gl_rom_n_890, ZN => gl_rom_n_1276);
  gl_rom_g35404 : ND4D0BWP7T port map(A1 => gl_rom_n_887, A2 => gl_rom_n_888, A3 => gl_rom_n_876, A4 => gl_rom_n_869, ZN => gl_rom_n_1275);
  gl_rom_g35405 : ND4D0BWP7T port map(A1 => gl_rom_n_882, A2 => gl_rom_n_886, A3 => gl_rom_n_883, A4 => gl_rom_n_884, ZN => gl_rom_n_1274);
  gl_rom_g35406 : ND4D0BWP7T port map(A1 => gl_rom_n_874, A2 => gl_rom_n_878, A3 => gl_rom_n_871, A4 => gl_rom_n_865, ZN => gl_rom_n_1273);
  gl_rom_g35407 : ND4D0BWP7T port map(A1 => gl_rom_n_873, A2 => gl_rom_n_881, A3 => gl_rom_n_875, A4 => gl_rom_n_877, ZN => gl_rom_n_1272);
  gl_rom_g35408 : ND4D0BWP7T port map(A1 => gl_rom_n_864, A2 => gl_rom_n_870, A3 => gl_rom_n_866, A4 => gl_rom_n_868, ZN => gl_rom_n_1271);
  gl_rom_g35409 : ND4D0BWP7T port map(A1 => gl_rom_n_862, A2 => gl_rom_n_856, A3 => gl_rom_n_854, A4 => gl_rom_n_859, ZN => gl_rom_n_1270);
  gl_rom_g35410 : ND4D0BWP7T port map(A1 => gl_rom_n_855, A2 => gl_rom_n_858, A3 => gl_rom_n_852, A4 => gl_rom_n_847, ZN => gl_rom_n_1269);
  gl_rom_g35411 : ND4D0BWP7T port map(A1 => gl_rom_n_848, A2 => gl_rom_n_853, A3 => gl_rom_n_849, A4 => gl_rom_n_851, ZN => gl_rom_n_1268);
  gl_rom_g35412 : ND4D0BWP7T port map(A1 => gl_rom_n_850, A2 => gl_rom_n_857, A3 => gl_rom_n_845, A4 => gl_rom_n_838, ZN => gl_rom_n_1267);
  gl_rom_g35413 : ND4D0BWP7T port map(A1 => gl_rom_n_846, A2 => gl_rom_n_841, A3 => gl_rom_n_843, A4 => gl_rom_n_840, ZN => gl_rom_n_1266);
  gl_rom_g35414 : ND4D0BWP7T port map(A1 => gl_rom_n_842, A2 => gl_rom_n_844, A3 => gl_rom_n_837, A4 => gl_rom_n_835, ZN => gl_rom_n_1265);
  gl_rom_g35415 : ND4D0BWP7T port map(A1 => gl_rom_n_872, A2 => gl_rom_n_755, A3 => gl_rom_n_706, A4 => gl_rom_n_816, ZN => gl_rom_n_1264);
  gl_rom_g35416 : ND4D0BWP7T port map(A1 => gl_rom_n_836, A2 => gl_rom_n_839, A3 => gl_rom_n_834, A4 => gl_rom_n_833, ZN => gl_rom_n_1263);
  gl_rom_g35417 : ND4D0BWP7T port map(A1 => gl_rom_n_798, A2 => gl_rom_n_824, A3 => gl_rom_n_767, A4 => gl_rom_n_742, ZN => gl_rom_n_1262);
  gl_rom_g35418 : ND4D0BWP7T port map(A1 => gl_rom_n_811, A2 => gl_rom_n_831, A3 => gl_rom_n_802, A4 => gl_rom_n_783, ZN => gl_rom_n_1261);
  gl_rom_g35419 : ND4D0BWP7T port map(A1 => gl_rom_n_826, A2 => gl_rom_n_832, A3 => gl_rom_n_828, A4 => gl_rom_n_830, ZN => gl_rom_n_1260);
  gl_rom_g35420 : ND4D0BWP7T port map(A1 => gl_rom_n_817, A2 => gl_rom_n_827, A3 => gl_rom_n_814, A4 => gl_rom_n_1062, ZN => gl_rom_n_1259);
  gl_rom_g35421 : ND4D0BWP7T port map(A1 => gl_rom_n_825, A2 => gl_rom_n_829, A3 => gl_rom_n_822, A4 => gl_rom_n_820, ZN => gl_rom_n_1258);
  gl_rom_g35422 : ND4D0BWP7T port map(A1 => gl_rom_n_818, A2 => gl_rom_n_823, A3 => gl_rom_n_819, A4 => gl_rom_n_821, ZN => gl_rom_n_1257);
  gl_rom_g35423 : ND4D0BWP7T port map(A1 => gl_rom_n_810, A2 => gl_rom_n_815, A3 => gl_rom_n_807, A4 => gl_rom_n_805, ZN => gl_rom_n_1256);
  gl_rom_g35424 : ND4D0BWP7T port map(A1 => gl_rom_n_809, A2 => gl_rom_n_813, A3 => gl_rom_n_812, A4 => gl_rom_n_808, ZN => gl_rom_n_1255);
  gl_rom_g35425 : ND4D0BWP7T port map(A1 => gl_rom_n_801, A2 => gl_rom_n_804, A3 => gl_rom_n_803, A4 => gl_rom_n_800, ZN => gl_rom_n_1254);
  gl_rom_g35426 : ND4D0BWP7T port map(A1 => gl_rom_n_791, A2 => gl_rom_n_797, A3 => gl_rom_n_782, A4 => gl_rom_n_778, ZN => gl_rom_n_1253);
  gl_rom_g35427 : ND4D0BWP7T port map(A1 => gl_rom_n_793, A2 => gl_rom_n_799, A3 => gl_rom_n_794, A4 => gl_rom_n_796, ZN => gl_rom_n_1252);
  gl_rom_g35428 : ND4D0BWP7T port map(A1 => gl_rom_n_792, A2 => gl_rom_n_795, A3 => gl_rom_n_788, A4 => gl_rom_n_785, ZN => gl_rom_n_1251);
  gl_rom_g35429 : ND4D0BWP7T port map(A1 => gl_rom_n_790, A2 => gl_rom_n_787, A3 => gl_rom_n_786, A4 => gl_rom_n_789, ZN => gl_rom_n_1250);
  gl_rom_g35430 : ND4D0BWP7T port map(A1 => gl_rom_n_781, A2 => gl_rom_n_776, A3 => gl_rom_n_769, A4 => gl_rom_n_774, ZN => gl_rom_n_1249);
  gl_rom_g35431 : ND4D0BWP7T port map(A1 => gl_rom_n_784, A2 => gl_rom_n_779, A3 => gl_rom_n_777, A4 => gl_rom_n_780, ZN => gl_rom_n_1248);
  gl_rom_g35432 : ND4D0BWP7T port map(A1 => gl_rom_n_775, A2 => gl_rom_n_772, A3 => gl_rom_n_773, A4 => gl_rom_n_768, ZN => gl_rom_n_1247);
  gl_rom_g35433 : ND4D0BWP7T port map(A1 => gl_rom_n_766, A2 => gl_rom_n_763, A3 => gl_rom_n_762, A4 => gl_rom_n_765, ZN => gl_rom_n_1246);
  gl_rom_g35434 : ND4D0BWP7T port map(A1 => gl_rom_n_760, A2 => gl_rom_n_770, A3 => gl_rom_n_741, A4 => gl_rom_n_734, ZN => gl_rom_n_1245);
  gl_rom_g35435 : ND4D0BWP7T port map(A1 => gl_rom_n_753, A2 => gl_rom_n_764, A3 => gl_rom_n_757, A4 => gl_rom_n_761, ZN => gl_rom_n_1244);
  gl_rom_g35436 : ND4D0BWP7T port map(A1 => gl_rom_n_759, A2 => gl_rom_n_743, A3 => gl_rom_n_731, A4 => gl_rom_n_751, ZN => gl_rom_n_1243);
  gl_rom_g35437 : ND4D0BWP7T port map(A1 => gl_rom_n_752, A2 => gl_rom_n_758, A3 => gl_rom_n_754, A4 => gl_rom_n_756, ZN => gl_rom_n_1242);
  gl_rom_g35438 : ND4D0BWP7T port map(A1 => gl_rom_n_749, A2 => gl_rom_n_745, A3 => gl_rom_n_744, A4 => gl_rom_n_747, ZN => gl_rom_n_1241);
  gl_rom_g35439 : ND4D0BWP7T port map(A1 => gl_rom_n_748, A2 => gl_rom_n_739, A3 => gl_rom_n_735, A4 => gl_rom_n_746, ZN => gl_rom_n_1240);
  gl_rom_g35440 : ND4D0BWP7T port map(A1 => gl_rom_n_738, A2 => gl_rom_n_740, A3 => gl_rom_n_737, A4 => gl_rom_n_736, ZN => gl_rom_n_1239);
  gl_rom_g35441 : ND4D0BWP7T port map(A1 => gl_rom_n_722, A2 => gl_rom_n_726, A3 => gl_rom_n_712, A4 => gl_rom_n_708, ZN => gl_rom_n_1238);
  gl_rom_g35442 : ND4D0BWP7T port map(A1 => gl_rom_n_733, A2 => gl_rom_n_729, A3 => gl_rom_n_728, A4 => gl_rom_n_732, ZN => gl_rom_n_1237);
  gl_rom_g35443 : ND4D0BWP7T port map(A1 => gl_rom_n_727, A2 => gl_rom_n_730, A3 => gl_rom_n_724, A4 => gl_rom_n_719, ZN => gl_rom_n_1236);
  gl_rom_g35444 : ND4D0BWP7T port map(A1 => gl_rom_n_725, A2 => gl_rom_n_721, A3 => gl_rom_n_723, A4 => gl_rom_n_720, ZN => gl_rom_n_1235);
  gl_rom_g35445 : ND4D0BWP7T port map(A1 => gl_rom_n_716, A2 => gl_rom_n_710, A3 => gl_rom_n_714, A4 => gl_rom_n_705, ZN => gl_rom_n_1234);
  gl_rom_g35446 : ND4D0BWP7T port map(A1 => gl_rom_n_718, A2 => gl_rom_n_715, A3 => gl_rom_n_713, A4 => gl_rom_n_717, ZN => gl_rom_n_1233);
  gl_rom_g35447 : ND4D0BWP7T port map(A1 => gl_rom_n_709, A2 => gl_rom_n_711, A3 => gl_rom_n_707, A4 => gl_rom_n_704, ZN => gl_rom_n_1232);
  gl_rom_g35448 : ND4D0BWP7T port map(A1 => gl_rom_n_703, A2 => gl_rom_n_698, A3 => gl_rom_n_636, A4 => gl_rom_n_639, ZN => gl_rom_n_1231);
  gl_rom_g35449 : ND4D0BWP7T port map(A1 => gl_rom_n_701, A2 => gl_rom_n_702, A3 => gl_rom_n_699, A4 => gl_rom_n_696, ZN => gl_rom_n_1230);
  gl_rom_g35450 : ND4D0BWP7T port map(A1 => gl_rom_n_700, A2 => gl_rom_n_691, A3 => gl_rom_n_697, A4 => gl_rom_n_688, ZN => gl_rom_n_1229);
  gl_rom_g35451 : ND4D0BWP7T port map(A1 => gl_rom_n_694, A2 => gl_rom_n_690, A3 => gl_rom_n_692, A4 => gl_rom_n_687, ZN => gl_rom_n_1228);
  gl_rom_g35452 : ND4D0BWP7T port map(A1 => gl_rom_n_695, A2 => gl_rom_n_683, A3 => gl_rom_n_672, A4 => gl_rom_n_689, ZN => gl_rom_n_1227);
  gl_rom_g35453 : ND4D0BWP7T port map(A1 => gl_rom_n_686, A2 => gl_rom_n_682, A3 => gl_rom_n_675, A4 => gl_rom_n_678, ZN => gl_rom_n_1226);
  gl_rom_g35454 : ND4D0BWP7T port map(A1 => gl_rom_n_680, A2 => gl_rom_n_685, A3 => gl_rom_n_681, A4 => gl_rom_n_684, ZN => gl_rom_n_1225);
  gl_rom_g35455 : ND4D0BWP7T port map(A1 => gl_rom_n_673, A2 => gl_rom_n_677, A3 => gl_rom_n_674, A4 => gl_rom_n_676, ZN => gl_rom_n_1224);
  gl_rom_g35456 : ND4D0BWP7T port map(A1 => gl_rom_n_679, A2 => gl_rom_n_693, A3 => gl_rom_n_669, A4 => gl_rom_n_652, ZN => gl_rom_n_1223);
  gl_rom_g35457 : ND4D0BWP7T port map(A1 => gl_rom_n_667, A2 => gl_rom_n_671, A3 => gl_rom_n_670, A4 => gl_rom_n_666, ZN => gl_rom_n_1222);
  gl_rom_g35458 : ND4D0BWP7T port map(A1 => gl_rom_n_668, A2 => gl_rom_n_660, A3 => gl_rom_n_657, A4 => gl_rom_n_664, ZN => gl_rom_n_1221);
  gl_rom_g35459 : ND4D0BWP7T port map(A1 => gl_rom_n_665, A2 => gl_rom_n_655, A3 => gl_rom_n_648, A4 => gl_rom_n_663, ZN => gl_rom_n_1220);
  gl_rom_g35460 : ND4D0BWP7T port map(A1 => gl_rom_n_662, A2 => gl_rom_n_661, A3 => gl_rom_n_658, A4 => gl_rom_n_659, ZN => gl_rom_n_1219);
  gl_rom_g35461 : ND4D0BWP7T port map(A1 => gl_rom_n_653, A2 => gl_rom_n_650, A3 => gl_rom_n_643, A4 => gl_rom_n_645, ZN => gl_rom_n_1218);
  gl_rom_g35462 : ND4D0BWP7T port map(A1 => gl_rom_n_649, A2 => gl_rom_n_656, A3 => gl_rom_n_651, A4 => gl_rom_n_654, ZN => gl_rom_n_1217);
  gl_rom_g35463 : ND4D0BWP7T port map(A1 => gl_rom_n_644, A2 => gl_rom_n_647, A3 => gl_rom_n_646, A4 => gl_rom_n_642, ZN => gl_rom_n_1216);
  gl_rom_g35464 : ND4D0BWP7T port map(A1 => gl_rom_n_634, A2 => gl_rom_n_640, A3 => gl_rom_n_635, A4 => gl_rom_n_638, ZN => gl_rom_n_1215);
  gl_rom_g35465 : ND4D0BWP7T port map(A1 => gl_rom_n_623, A2 => gl_rom_n_628, A3 => gl_rom_n_608, A4 => gl_rom_n_589, ZN => gl_rom_n_1214);
  gl_rom_g35466 : ND4D0BWP7T port map(A1 => gl_rom_n_637, A2 => gl_rom_n_630, A3 => gl_rom_n_627, A4 => gl_rom_n_633, ZN => gl_rom_n_1213);
  gl_rom_g35467 : ND4D0BWP7T port map(A1 => gl_rom_n_632, A2 => gl_rom_n_619, A3 => gl_rom_n_616, A4 => gl_rom_n_624, ZN => gl_rom_n_1212);
  gl_rom_g35468 : ND4D0BWP7T port map(A1 => gl_rom_n_626, A2 => gl_rom_n_631, A3 => gl_rom_n_629, A4 => gl_rom_n_625, ZN => gl_rom_n_1211);
  gl_rom_g35469 : ND4D0BWP7T port map(A1 => gl_rom_n_615, A2 => gl_rom_n_622, A3 => gl_rom_n_617, A4 => gl_rom_n_620, ZN => gl_rom_n_1210);
  gl_rom_g35470 : ND4D0BWP7T port map(A1 => gl_rom_n_609, A2 => gl_rom_n_621, A3 => gl_rom_n_614, A4 => gl_rom_n_618, ZN => gl_rom_n_1209);
  gl_rom_g35471 : ND4D0BWP7T port map(A1 => gl_rom_n_610, A2 => gl_rom_n_613, A3 => gl_rom_n_611, A4 => gl_rom_n_612, ZN => gl_rom_n_1208);
  gl_rom_g35472 : ND4D0BWP7T port map(A1 => gl_rom_n_600, A2 => gl_rom_n_588, A3 => gl_rom_n_581, A4 => gl_rom_n_596, ZN => gl_rom_n_1207);
  gl_rom_g35473 : ND4D0BWP7T port map(A1 => gl_rom_n_606, A2 => gl_rom_n_607, A3 => gl_rom_n_603, A4 => gl_rom_n_602, ZN => gl_rom_n_1206);
  gl_rom_g35474 : ND4D0BWP7T port map(A1 => gl_rom_n_601, A2 => gl_rom_n_605, A3 => gl_rom_n_598, A4 => gl_rom_n_593, ZN => gl_rom_n_1205);
  gl_rom_g35475 : ND4D0BWP7T port map(A1 => gl_rom_n_599, A2 => gl_rom_n_595, A3 => gl_rom_n_594, A4 => gl_rom_n_597, ZN => gl_rom_n_1204);
  gl_rom_g35476 : ND4D0BWP7T port map(A1 => gl_rom_n_591, A2 => gl_rom_n_585, A3 => gl_rom_n_579, A4 => gl_rom_n_584, ZN => gl_rom_n_1203);
  gl_rom_g35477 : ND4D0BWP7T port map(A1 => gl_rom_n_586, A2 => gl_rom_n_592, A3 => gl_rom_n_587, A4 => gl_rom_n_590, ZN => gl_rom_n_1202);
  gl_rom_g35478 : ND4D0BWP7T port map(A1 => gl_rom_n_583, A2 => gl_rom_n_580, A3 => gl_rom_n_578, A4 => gl_rom_n_582, ZN => gl_rom_n_1201);
  gl_rom_g35479 : ND4D0BWP7T port map(A1 => gl_rom_n_604, A2 => gl_rom_n_577, A3 => gl_rom_n_455, A4 => gl_rom_n_482, ZN => gl_rom_n_1200);
  gl_rom_g35480 : ND4D0BWP7T port map(A1 => gl_rom_n_545, A2 => gl_rom_n_575, A3 => gl_rom_n_514, A4 => gl_rom_n_490, ZN => gl_rom_n_1199);
  gl_rom_g35481 : ND4D0BWP7T port map(A1 => gl_rom_n_569, A2 => gl_rom_n_576, A3 => gl_rom_n_572, A4 => gl_rom_n_573, ZN => gl_rom_n_1198);
  gl_rom_g35482 : ND4D0BWP7T port map(A1 => gl_rom_n_558, A2 => gl_rom_n_568, A3 => gl_rom_n_542, A4 => gl_rom_n_529, ZN => gl_rom_n_1197);
  gl_rom_g35483 : ND4D0BWP7T port map(A1 => gl_rom_n_574, A2 => gl_rom_n_570, A3 => gl_rom_n_564, A4 => gl_rom_n_566, ZN => gl_rom_n_1196);
  gl_rom_g35484 : ND4D0BWP7T port map(A1 => gl_rom_n_571, A2 => gl_rom_n_554, A3 => gl_rom_n_551, A4 => gl_rom_n_561, ZN => gl_rom_n_1195);
  gl_rom_g35485 : ND4D0BWP7T port map(A1 => gl_rom_n_567, A2 => gl_rom_n_563, A3 => gl_rom_n_562, A4 => gl_rom_n_565, ZN => gl_rom_n_1194);
  gl_rom_g35486 : ND4D0BWP7T port map(A1 => gl_rom_n_556, A2 => gl_rom_n_560, A3 => gl_rom_n_552, A4 => gl_rom_n_548, ZN => gl_rom_n_1193);
  gl_rom_g35487 : ND4D0BWP7T port map(A1 => gl_rom_n_553, A2 => gl_rom_n_559, A3 => gl_rom_n_555, A4 => gl_rom_n_557, ZN => gl_rom_n_1192);
  gl_rom_g35488 : ND4D0BWP7T port map(A1 => gl_rom_n_641, A2 => gl_rom_n_910, A3 => gl_rom_n_750, A4 => gl_rom_n_861, ZN => gl_rom_n_1191);
  gl_rom_g35489 : ND4D0BWP7T port map(A1 => gl_rom_n_44, A2 => gl_rom_n_41, A3 => gl_rom_n_806, A4 => gl_rom_n_39, ZN => gl_rom_n_1190);
  gl_rom_g35490 : ND4D0BWP7T port map(A1 => gl_rom_n_537, A2 => gl_rom_n_544, A3 => gl_rom_n_539, A4 => gl_rom_n_543, ZN => gl_rom_n_1189);
  gl_rom_g35491 : ND4D0BWP7T port map(A1 => gl_rom_n_541, A2 => gl_rom_n_535, A3 => gl_rom_n_531, A4 => gl_rom_n_538, ZN => gl_rom_n_1188);
  gl_rom_g35492 : ND4D0BWP7T port map(A1 => gl_rom_n_530, A2 => gl_rom_n_536, A3 => gl_rom_n_532, A4 => gl_rom_n_534, ZN => gl_rom_n_1187);
  gl_rom_g35493 : ND4D0BWP7T port map(A1 => gl_rom_n_526, A2 => gl_rom_n_528, A3 => gl_rom_n_523, A4 => gl_rom_n_522, ZN => gl_rom_n_1186);
  gl_rom_g35494 : ND4D0BWP7T port map(A1 => gl_rom_n_524, A2 => gl_rom_n_525, A3 => gl_rom_n_519, A4 => gl_rom_n_517, ZN => gl_rom_n_1185);
  gl_rom_g35495 : ND4D0BWP7T port map(A1 => gl_rom_n_518, A2 => gl_rom_n_521, A3 => gl_rom_n_516, A4 => gl_rom_n_515, ZN => gl_rom_n_1184);
  gl_rom_g35496 : ND4D0BWP7T port map(A1 => gl_rom_n_498, A2 => gl_rom_n_510, A3 => gl_rom_n_480, A4 => gl_rom_n_476, ZN => gl_rom_n_1183);
  gl_rom_g35497 : ND4D0BWP7T port map(A1 => gl_rom_n_513, A2 => gl_rom_n_509, A3 => gl_rom_n_508, A4 => gl_rom_n_512, ZN => gl_rom_n_1182);
  gl_rom_g35498 : ND4D0BWP7T port map(A1 => gl_rom_n_504, A2 => gl_rom_n_511, A3 => gl_rom_n_507, A4 => gl_rom_n_501, ZN => gl_rom_n_1181);
  gl_rom_g35499 : ND4D0BWP7T port map(A1 => gl_rom_n_505, A2 => gl_rom_n_493, A3 => gl_rom_n_487, A4 => gl_rom_n_502, ZN => gl_rom_n_1180);
  gl_rom_g35500 : ND4D0BWP7T port map(A1 => gl_rom_n_503, A2 => gl_rom_n_506, A3 => gl_rom_n_500, A4 => gl_rom_n_499, ZN => gl_rom_n_1179);
  gl_rom_g35501 : ND4D0BWP7T port map(A1 => gl_rom_n_425, A2 => gl_rom_n_271, A3 => gl_rom_n_203, A4 => gl_rom_n_326, ZN => gl_rom_n_1178);
  gl_rom_g35502 : ND4D0BWP7T port map(A1 => gl_rom_n_485, A2 => gl_rom_n_496, A3 => gl_rom_n_488, A4 => gl_rom_n_492, ZN => gl_rom_n_1177);
  gl_rom_g35503 : ND4D0BWP7T port map(A1 => gl_rom_n_491, A2 => gl_rom_n_497, A3 => gl_rom_n_494, A4 => gl_rom_n_495, ZN => gl_rom_n_1176);
  gl_rom_g35504 : ND4D0BWP7T port map(A1 => gl_rom_n_483, A2 => gl_rom_n_489, A3 => gl_rom_n_484, A4 => gl_rom_n_486, ZN => gl_rom_n_1175);
  gl_rom_g35505 : ND4D0BWP7T port map(A1 => gl_rom_n_474, A2 => gl_rom_n_481, A3 => gl_rom_n_477, A4 => gl_rom_n_479, ZN => gl_rom_n_1174);
  gl_rom_g35506 : ND4D0BWP7T port map(A1 => gl_rom_n_475, A2 => gl_rom_n_478, A3 => gl_rom_n_469, A4 => gl_rom_n_467, ZN => gl_rom_n_1173);
  gl_rom_g35507 : ND4D0BWP7T port map(A1 => gl_rom_n_473, A2 => gl_rom_n_462, A3 => gl_rom_n_454, A4 => gl_rom_n_471, ZN => gl_rom_n_1172);
  gl_rom_g35508 : ND4D0BWP7T port map(A1 => gl_rom_n_466, A2 => gl_rom_n_472, A3 => gl_rom_n_468, A4 => gl_rom_n_470, ZN => gl_rom_n_1171);
  gl_rom_g35509 : ND4D0BWP7T port map(A1 => gl_rom_n_419, A2 => gl_rom_n_450, A3 => gl_rom_n_386, A4 => gl_rom_n_363, ZN => gl_rom_n_1170);
  gl_rom_g35510 : ND4D0BWP7T port map(A1 => gl_rom_n_464, A2 => gl_rom_n_457, A3 => gl_rom_n_452, A4 => gl_rom_n_460, ZN => gl_rom_n_1169);
  gl_rom_g35511 : ND4D0BWP7T port map(A1 => gl_rom_n_465, A2 => gl_rom_n_461, A3 => gl_rom_n_459, A4 => gl_rom_n_463, ZN => gl_rom_n_1168);
  gl_rom_g35512 : ND4D0BWP7T port map(A1 => gl_rom_n_458, A2 => gl_rom_n_453, A3 => gl_rom_n_451, A4 => gl_rom_n_456, ZN => gl_rom_n_1167);
  gl_rom_g35513 : ND4D0BWP7T port map(A1 => gl_rom_n_449, A2 => gl_rom_n_446, A3 => gl_rom_n_443, A4 => gl_rom_n_447, ZN => gl_rom_n_1166);
  gl_rom_g35514 : ND4D0BWP7T port map(A1 => gl_rom_n_432, A2 => gl_rom_n_445, A3 => gl_rom_n_416, A4 => gl_rom_n_401, ZN => gl_rom_n_1165);
  gl_rom_g35515 : ND4D0BWP7T port map(A1 => gl_rom_n_448, A2 => gl_rom_n_440, A3 => gl_rom_n_438, A4 => gl_rom_n_444, ZN => gl_rom_n_1164);
  gl_rom_g35516 : ND4D0BWP7T port map(A1 => gl_rom_n_435, A2 => gl_rom_n_442, A3 => gl_rom_n_428, A4 => gl_rom_n_424, ZN => gl_rom_n_1163);
  gl_rom_g35517 : ND4D0BWP7T port map(A1 => gl_rom_n_436, A2 => gl_rom_n_441, A3 => gl_rom_n_437, A4 => gl_rom_n_439, ZN => gl_rom_n_1162);
  gl_rom_g35518 : ND4D0BWP7T port map(A1 => gl_rom_n_426, A2 => gl_rom_n_434, A3 => gl_rom_n_430, A4 => gl_rom_n_421, ZN => gl_rom_n_1161);
  gl_rom_g35519 : ND4D0BWP7T port map(A1 => gl_rom_n_427, A2 => gl_rom_n_433, A3 => gl_rom_n_429, A4 => gl_rom_n_431, ZN => gl_rom_n_1160);
  gl_rom_g35520 : ND4D0BWP7T port map(A1 => gl_rom_n_418, A2 => gl_rom_n_423, A3 => gl_rom_n_420, A4 => gl_rom_n_422, ZN => gl_rom_n_1159);
  gl_rom_g35521 : ND4D0BWP7T port map(A1 => gl_rom_n_417, A2 => gl_rom_n_413, A3 => gl_rom_n_411, A4 => gl_rom_n_415, ZN => gl_rom_n_1158);
  gl_rom_g35522 : ND4D0BWP7T port map(A1 => gl_rom_n_410, A2 => gl_rom_n_414, A3 => gl_rom_n_407, A4 => gl_rom_n_406, ZN => gl_rom_n_1157);
  gl_rom_g35523 : ND4D0BWP7T port map(A1 => gl_rom_n_403, A2 => gl_rom_n_412, A3 => gl_rom_n_398, A4 => gl_rom_n_393, ZN => gl_rom_n_1156);
  gl_rom_g35524 : ND4D0BWP7T port map(A1 => gl_rom_n_405, A2 => gl_rom_n_409, A3 => gl_rom_n_408, A4 => gl_rom_n_404, ZN => gl_rom_n_1155);
  gl_rom_g35525 : ND4D0BWP7T port map(A1 => gl_rom_n_395, A2 => gl_rom_n_402, A3 => gl_rom_n_397, A4 => gl_rom_n_399, ZN => gl_rom_n_1154);
  gl_rom_g35526 : ND4D0BWP7T port map(A1 => gl_rom_n_396, A2 => gl_rom_n_400, A3 => gl_rom_n_392, A4 => gl_rom_n_390, ZN => gl_rom_n_1153);
  gl_rom_g35527 : ND4D0BWP7T port map(A1 => gl_rom_n_388, A2 => gl_rom_n_394, A3 => gl_rom_n_389, A4 => gl_rom_n_391, ZN => gl_rom_n_1152);
  gl_rom_g35528 : ND4D0BWP7T port map(A1 => gl_rom_n_370, A2 => gl_rom_n_384, A3 => gl_rom_n_353, A4 => gl_rom_n_342, ZN => gl_rom_n_1151);
  gl_rom_g35529 : ND4D0BWP7T port map(A1 => gl_rom_n_379, A2 => gl_rom_n_385, A3 => gl_rom_n_381, A4 => gl_rom_n_383, ZN => gl_rom_n_1150);
  gl_rom_g35530 : ND4D0BWP7T port map(A1 => gl_rom_n_380, A2 => gl_rom_n_382, A3 => gl_rom_n_376, A4 => gl_rom_n_373, ZN => gl_rom_n_1149);
  gl_rom_g35531 : ND4D0BWP7T port map(A1 => gl_rom_n_378, A2 => gl_rom_n_362, A3 => gl_rom_n_359, A4 => gl_rom_n_374, ZN => gl_rom_n_1148);
  gl_rom_g35532 : ND4D0BWP7T port map(A1 => gl_rom_n_371, A2 => gl_rom_n_377, A3 => gl_rom_n_372, A4 => gl_rom_n_375, ZN => gl_rom_n_1147);
  gl_rom_g35533 : ND4D0BWP7T port map(A1 => gl_rom_n_368, A2 => gl_rom_n_361, A3 => gl_rom_n_357, A4 => gl_rom_n_365, ZN => gl_rom_n_1146);
  gl_rom_g35534 : ND4D0BWP7T port map(A1 => gl_rom_n_367, A2 => gl_rom_n_369, A3 => gl_rom_n_366, A4 => gl_rom_n_364, ZN => gl_rom_n_1145);
  gl_rom_g35535 : ND4D0BWP7T port map(A1 => gl_rom_n_360, A2 => gl_rom_n_358, A3 => gl_rom_n_355, A4 => gl_rom_n_356, ZN => gl_rom_n_1144);
  gl_rom_g35536 : ND4D0BWP7T port map(A1 => gl_rom_n_350, A2 => gl_rom_n_331, A3 => gl_rom_n_329, A4 => gl_rom_n_341, ZN => gl_rom_n_1143);
  gl_rom_g35537 : ND4D0BWP7T port map(A1 => gl_rom_n_354, A2 => gl_rom_n_349, A3 => gl_rom_n_347, A4 => gl_rom_n_351, ZN => gl_rom_n_1142);
  gl_rom_g35538 : ND4D0BWP7T port map(A1 => gl_rom_n_348, A2 => gl_rom_n_352, A3 => gl_rom_n_343, A4 => gl_rom_n_339, ZN => gl_rom_n_1141);
  gl_rom_g35539 : ND4D0BWP7T port map(A1 => gl_rom_n_346, A2 => gl_rom_n_340, A3 => gl_rom_n_338, A4 => gl_rom_n_344, ZN => gl_rom_n_1140);
  gl_rom_g35540 : ND4D0BWP7T port map(A1 => gl_rom_n_345, A2 => gl_rom_n_289, A3 => gl_rom_n_257, A4 => gl_rom_n_265, ZN => gl_rom_n_1139);
  gl_rom_g35541 : ND4D0BWP7T port map(A1 => gl_rom_n_336, A2 => gl_rom_n_328, A3 => gl_rom_n_325, A4 => gl_rom_n_334, ZN => gl_rom_n_1138);
  gl_rom_g35542 : ND4D0BWP7T port map(A1 => gl_rom_n_332, A2 => gl_rom_n_337, A3 => gl_rom_n_333, A4 => gl_rom_n_335, ZN => gl_rom_n_1137);
  gl_rom_g35543 : ND4D0BWP7T port map(A1 => gl_rom_n_323, A2 => gl_rom_n_330, A3 => gl_rom_n_324, A4 => gl_rom_n_327, ZN => gl_rom_n_1136);
  gl_rom_g35544 : ND4D0BWP7T port map(A1 => gl_rom_n_302, A2 => gl_rom_n_322, A3 => gl_rom_n_288, A4 => gl_rom_n_279, ZN => gl_rom_n_1135);
  gl_rom_g35545 : ND4D0BWP7T port map(A1 => gl_rom_n_321, A2 => gl_rom_n_318, A3 => gl_rom_n_315, A4 => gl_rom_n_319, ZN => gl_rom_n_1134);
  gl_rom_g35546 : ND4D0BWP7T port map(A1 => gl_rom_n_317, A2 => gl_rom_n_298, A3 => gl_rom_n_293, A4 => gl_rom_n_309, ZN => gl_rom_n_1133);
  gl_rom_g35547 : ND4D0BWP7T port map(A1 => gl_rom_n_316, A2 => gl_rom_n_320, A3 => gl_rom_n_312, A4 => gl_rom_n_308, ZN => gl_rom_n_1132);
  gl_rom_g35548 : ND4D0BWP7T port map(A1 => gl_rom_n_313, A2 => gl_rom_n_314, A3 => gl_rom_n_304, A4 => gl_rom_n_301, ZN => gl_rom_n_1131);
  gl_rom_g35549 : ND4D0BWP7T port map(A1 => gl_rom_n_306, A2 => gl_rom_n_311, A3 => gl_rom_n_307, A4 => gl_rom_n_310, ZN => gl_rom_n_1130);
  gl_rom_g35550 : ND4D0BWP7T port map(A1 => gl_rom_n_303, A2 => gl_rom_n_305, A3 => gl_rom_n_300, A4 => gl_rom_n_299, ZN => gl_rom_n_1129);
  gl_rom_g35551 : ND4D0BWP7T port map(A1 => gl_rom_n_297, A2 => gl_rom_n_291, A3 => gl_rom_n_286, A4 => gl_rom_n_296, ZN => gl_rom_n_1128);
  gl_rom_g35552 : ND4D0BWP7T port map(A1 => gl_rom_n_290, A2 => gl_rom_n_295, A3 => gl_rom_n_292, A4 => gl_rom_n_550, ZN => gl_rom_n_1127);
  gl_rom_g35553 : ND4D0BWP7T port map(A1 => gl_rom_n_285, A2 => gl_rom_n_287, A3 => gl_rom_n_284, A4 => gl_rom_n_283, ZN => gl_rom_n_1126);
  gl_rom_g35554 : ND4D0BWP7T port map(A1 => gl_rom_n_281, A2 => gl_rom_n_282, A3 => gl_rom_n_270, A4 => gl_rom_n_262, ZN => gl_rom_n_1125);
  gl_rom_g35555 : ND4D0BWP7T port map(A1 => gl_rom_n_274, A2 => gl_rom_n_280, A3 => gl_rom_n_276, A4 => gl_rom_n_278, ZN => gl_rom_n_1124);
  gl_rom_g35556 : ND4D0BWP7T port map(A1 => gl_rom_n_266, A2 => gl_rom_n_277, A3 => gl_rom_n_269, A4 => gl_rom_n_275, ZN => gl_rom_n_1123);
  gl_rom_g35557 : ND4D0BWP7T port map(A1 => gl_rom_n_272, A2 => gl_rom_n_273, A3 => gl_rom_n_268, A4 => gl_rom_n_267, ZN => gl_rom_n_1122);
  gl_rom_g35558 : ND4D0BWP7T port map(A1 => gl_rom_n_261, A2 => gl_rom_n_254, A3 => gl_rom_n_251, A4 => gl_rom_n_259, ZN => gl_rom_n_1121);
  gl_rom_g35559 : ND4D0BWP7T port map(A1 => gl_rom_n_258, A2 => gl_rom_n_264, A3 => gl_rom_n_260, A4 => gl_rom_n_263, ZN => gl_rom_n_1120);
  gl_rom_g35560 : ND4D0BWP7T port map(A1 => gl_rom_n_256, A2 => gl_rom_n_252, A3 => gl_rom_n_255, A4 => gl_rom_n_250, ZN => gl_rom_n_1119);
  gl_rom_g35561 : ND4D0BWP7T port map(A1 => gl_rom_n_249, A2 => gl_rom_n_253, A3 => gl_rom_n_231, A4 => gl_rom_n_219, ZN => gl_rom_n_1118);
  gl_rom_g35562 : ND4D0BWP7T port map(A1 => gl_rom_n_248, A2 => gl_rom_n_245, A3 => gl_rom_n_247, A4 => gl_rom_n_244, ZN => gl_rom_n_1117);
  gl_rom_g35563 : ND4D0BWP7T port map(A1 => gl_rom_n_243, A2 => gl_rom_n_246, A3 => gl_rom_n_238, A4 => gl_rom_n_236, ZN => gl_rom_n_1116);
  gl_rom_g35564 : ND4D0BWP7T port map(A1 => gl_rom_n_240, A2 => gl_rom_n_242, A3 => gl_rom_n_230, A4 => gl_rom_n_226, ZN => gl_rom_n_1115);
  gl_rom_g35565 : ND4D0BWP7T port map(A1 => gl_rom_n_239, A2 => gl_rom_n_241, A3 => gl_rom_n_237, A4 => gl_rom_n_235, ZN => gl_rom_n_1114);
  gl_rom_g35566 : ND4D0BWP7T port map(A1 => gl_rom_n_227, A2 => gl_rom_n_232, A3 => gl_rom_n_224, A4 => gl_rom_n_222, ZN => gl_rom_n_1113);
  gl_rom_g35567 : ND4D0BWP7T port map(A1 => gl_rom_n_234, A2 => gl_rom_n_229, A3 => gl_rom_n_228, A4 => gl_rom_n_233, ZN => gl_rom_n_1112);
  gl_rom_g35568 : ND4D0BWP7T port map(A1 => gl_rom_n_221, A2 => gl_rom_n_225, A3 => gl_rom_n_223, A4 => gl_rom_n_220, ZN => gl_rom_n_1111);
  gl_rom_g35569 : ND4D0BWP7T port map(A1 => gl_rom_n_218, A2 => gl_rom_n_215, A3 => gl_rom_n_214, A4 => gl_rom_n_217, ZN => gl_rom_n_1110);
  gl_rom_g35570 : ND4D0BWP7T port map(A1 => gl_rom_n_191, A2 => gl_rom_n_172, A3 => gl_rom_n_116, A4 => gl_rom_n_144, ZN => gl_rom_n_1109);
  gl_rom_g35571 : ND4D0BWP7T port map(A1 => gl_rom_n_216, A2 => gl_rom_n_208, A3 => gl_rom_n_205, A4 => gl_rom_n_212, ZN => gl_rom_n_1108);
  gl_rom_g35572 : ND4D0BWP7T port map(A1 => gl_rom_n_211, A2 => gl_rom_n_213, A3 => gl_rom_n_202, A4 => gl_rom_n_194, ZN => gl_rom_n_1107);
  gl_rom_g35573 : ND4D0BWP7T port map(A1 => gl_rom_n_206, A2 => gl_rom_n_210, A3 => gl_rom_n_207, A4 => gl_rom_n_209, ZN => gl_rom_n_1106);
  gl_rom_g35574 : ND4D0BWP7T port map(A1 => gl_rom_n_198, A2 => gl_rom_n_200, A3 => gl_rom_n_193, A4 => gl_rom_n_189, ZN => gl_rom_n_1105);
  gl_rom_g35575 : ND4D0BWP7T port map(A1 => gl_rom_n_204, A2 => gl_rom_n_199, A3 => gl_rom_n_197, A4 => gl_rom_n_201, ZN => gl_rom_n_1104);
  gl_rom_g35576 : ND4D0BWP7T port map(A1 => gl_rom_n_192, A2 => gl_rom_n_195, A3 => gl_rom_n_190, A4 => gl_rom_n_188, ZN => gl_rom_n_1103);
  gl_rom_g35577 : ND4D0BWP7T port map(A1 => gl_rom_n_187, A2 => gl_rom_n_186, A3 => gl_rom_n_182, A4 => gl_rom_n_184, ZN => gl_rom_n_1102);
  gl_rom_g35578 : ND4D0BWP7T port map(A1 => gl_rom_n_171, A2 => gl_rom_n_180, A3 => gl_rom_n_155, A4 => gl_rom_n_140, ZN => gl_rom_n_1101);
  gl_rom_g35579 : ND4D0BWP7T port map(A1 => gl_rom_n_181, A2 => gl_rom_n_185, A3 => gl_rom_n_177, A4 => gl_rom_n_175, ZN => gl_rom_n_1100);
  gl_rom_g35580 : ND4D0BWP7T port map(A1 => gl_rom_n_183, A2 => gl_rom_n_173, A3 => gl_rom_n_163, A4 => gl_rom_n_167, ZN => gl_rom_n_1099);
  gl_rom_g35581 : ND4D0BWP7T port map(A1 => gl_rom_n_179, A2 => gl_rom_n_178, A3 => gl_rom_n_174, A4 => gl_rom_n_176, ZN => gl_rom_n_1098);
  gl_rom_g35582 : ND4D0BWP7T port map(A1 => gl_rom_n_164, A2 => gl_rom_n_170, A3 => gl_rom_n_165, A4 => gl_rom_n_168, ZN => gl_rom_n_1097);
  gl_rom_g35583 : ND4D0BWP7T port map(A1 => gl_rom_n_169, A2 => gl_rom_n_162, A3 => gl_rom_n_166, A4 => gl_rom_n_157, ZN => gl_rom_n_1096);
  gl_rom_g35584 : ND4D0BWP7T port map(A1 => gl_rom_n_158, A2 => gl_rom_n_161, A3 => gl_rom_n_159, A4 => gl_rom_n_160, ZN => gl_rom_n_1095);
  gl_rom_g35585 : ND4D0BWP7T port map(A1 => gl_rom_n_146, A2 => gl_rom_n_153, A3 => gl_rom_n_137, A4 => gl_rom_n_132, ZN => gl_rom_n_1094);
  gl_rom_g35586 : ND4D0BWP7T port map(A1 => gl_rom_n_156, A2 => gl_rom_n_151, A3 => gl_rom_n_154, A4 => gl_rom_n_149, ZN => gl_rom_n_1093);
  gl_rom_g35587 : ND4D0BWP7T port map(A1 => gl_rom_n_150, A2 => gl_rom_n_152, A3 => gl_rom_n_145, A4 => gl_rom_n_141, ZN => gl_rom_n_1092);
  gl_rom_g35588 : ND4D0BWP7T port map(A1 => gl_rom_n_142, A2 => gl_rom_n_148, A3 => gl_rom_n_143, A4 => gl_rom_n_147, ZN => gl_rom_n_1091);
  gl_rom_g35589 : ND4D0BWP7T port map(A1 => gl_rom_n_136, A2 => gl_rom_n_130, A3 => gl_rom_n_127, A4 => gl_rom_n_134, ZN => gl_rom_n_1090);
  gl_rom_g35590 : ND4D0BWP7T port map(A1 => gl_rom_n_133, A2 => gl_rom_n_139, A3 => gl_rom_n_135, A4 => gl_rom_n_138, ZN => gl_rom_n_1089);
  gl_rom_g35591 : ND4D0BWP7T port map(A1 => gl_rom_n_126, A2 => gl_rom_n_131, A3 => gl_rom_n_128, A4 => gl_rom_n_129, ZN => gl_rom_n_1088);
  gl_rom_g35592 : ND4D0BWP7T port map(A1 => gl_rom_n_125, A2 => gl_rom_n_121, A3 => gl_rom_n_120, A4 => gl_rom_n_124, ZN => gl_rom_n_1087);
  gl_rom_g35593 : ND4D0BWP7T port map(A1 => gl_rom_n_72, A2 => gl_rom_n_94, A3 => gl_rom_n_1026, A4 => gl_rom_n_966, ZN => gl_rom_n_1086);
  gl_rom_g35594 : ND4D0BWP7T port map(A1 => gl_rom_n_109, A2 => gl_rom_n_119, A3 => gl_rom_n_92, A4 => gl_rom_n_76, ZN => gl_rom_n_1085);
  gl_rom_g35595 : ND4D0BWP7T port map(A1 => gl_rom_n_196, A2 => gl_rom_n_78, A3 => gl_rom_n_387, A4 => gl_rom_n_771, ZN => gl_rom_n_1084);
  gl_rom_g35596 : ND4D0BWP7T port map(A1 => gl_rom_n_123, A2 => gl_rom_n_113, A3 => gl_rom_n_112, A4 => gl_rom_n_118, ZN => gl_rom_n_1083);
  gl_rom_g35597 : ND4D0BWP7T port map(A1 => gl_rom_n_122, A2 => gl_rom_n_105, A3 => gl_rom_n_101, A4 => gl_rom_n_114, ZN => gl_rom_n_1082);
  gl_rom_g35598 : ND4D0BWP7T port map(A1 => gl_rom_n_110, A2 => gl_rom_n_117, A3 => gl_rom_n_111, A4 => gl_rom_n_115, ZN => gl_rom_n_1081);
  gl_rom_g35599 : ND4D0BWP7T port map(A1 => gl_rom_n_97, A2 => gl_rom_n_107, A3 => gl_rom_n_99, A4 => gl_rom_n_102, ZN => gl_rom_n_1080);
  gl_rom_g35600 : ND4D0BWP7T port map(A1 => gl_rom_n_103, A2 => gl_rom_n_108, A3 => gl_rom_n_104, A4 => gl_rom_n_106, ZN => gl_rom_n_1079);
  gl_rom_g35601 : ND4D0BWP7T port map(A1 => gl_rom_n_95, A2 => gl_rom_n_100, A3 => gl_rom_n_96, A4 => gl_rom_n_98, ZN => gl_rom_n_1078);
  gl_rom_g35602 : ND4D0BWP7T port map(A1 => gl_rom_n_93, A2 => gl_rom_n_88, A3 => gl_rom_n_87, A4 => gl_rom_n_91, ZN => gl_rom_n_1077);
  gl_rom_g35603 : ND4D0BWP7T port map(A1 => gl_rom_n_89, A2 => gl_rom_n_75, A3 => gl_rom_n_85, A4 => gl_rom_n_68, ZN => gl_rom_n_1076);
  gl_rom_g35604 : ND4D0BWP7T port map(A1 => gl_rom_n_86, A2 => gl_rom_n_90, A3 => gl_rom_n_82, A4 => gl_rom_n_79, ZN => gl_rom_n_1075);
  gl_rom_g35605 : ND4D0BWP7T port map(A1 => gl_rom_n_84, A2 => gl_rom_n_81, A3 => gl_rom_n_80, A4 => gl_rom_n_83, ZN => gl_rom_n_1074);
  gl_rom_g35606 : ND4D0BWP7T port map(A1 => gl_rom_n_70, A2 => gl_rom_n_73, A3 => gl_rom_n_65, A4 => gl_rom_n_63, ZN => gl_rom_n_1073);
  gl_rom_g35607 : ND4D0BWP7T port map(A1 => gl_rom_n_71, A2 => gl_rom_n_77, A3 => gl_rom_n_74, A4 => gl_rom_n_69, ZN => gl_rom_n_1072);
  gl_rom_g35608 : ND4D0BWP7T port map(A1 => gl_rom_n_62, A2 => gl_rom_n_67, A3 => gl_rom_n_64, A4 => gl_rom_n_66, ZN => gl_rom_n_1071);
  gl_rom_g35609 : ND4D0BWP7T port map(A1 => gl_rom_n_45, A2 => gl_rom_n_58, A3 => gl_rom_n_1053, A4 => gl_rom_n_1036, ZN => gl_rom_n_1070);
  gl_rom_g35610 : ND4D0BWP7T port map(A1 => gl_rom_n_61, A2 => gl_rom_n_56, A3 => gl_rom_n_60, A4 => gl_rom_n_54, ZN => gl_rom_n_1069);
  gl_rom_g35611 : ND4D0BWP7T port map(A1 => gl_rom_n_59, A2 => gl_rom_n_52, A3 => gl_rom_n_47, A4 => gl_rom_n_55, ZN => gl_rom_n_1068);
  gl_rom_g35612 : ND4D0BWP7T port map(A1 => gl_rom_n_50, A2 => gl_rom_n_57, A3 => gl_rom_n_43, A4 => gl_rom_n_1061, ZN => gl_rom_n_1067);
  gl_rom_g35613 : ND4D0BWP7T port map(A1 => gl_rom_n_53, A2 => gl_rom_n_49, A3 => gl_rom_n_48, A4 => gl_rom_n_51, ZN => gl_rom_n_1066);
  gl_rom_g35614 : ND4D0BWP7T port map(A1 => gl_rom_n_1055, A2 => gl_rom_n_46, A3 => gl_rom_n_1022, A4 => gl_rom_n_1004, ZN => gl_rom_n_1065);
  gl_rom_g35615 : ND4D0BWP7T port map(A1 => gl_rom_n_40, A2 => gl_rom_n_42, A3 => gl_rom_n_1060, A4 => gl_rom_n_1057, ZN => gl_rom_n_1064);
  gl_rom_g35616 : ND4D0BWP7T port map(A1 => gl_rom_n_540, A2 => gl_rom_n_527, A3 => gl_rom_n_520, A4 => gl_rom_n_533, ZN => gl_rom_n_1063);
  gl_rom_g35617 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_584(0), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_587(0), ZN => gl_rom_n_1062);
  gl_rom_g35618 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_840(0), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_843(0), ZN => gl_rom_n_1061);
  gl_rom_g35619 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_257(0), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_261(0), ZN => gl_rom_n_1060);
  gl_rom_g35620 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_1002(1), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_1007(1), ZN => gl_rom_n_1059);
  gl_rom_g35621 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_1001(1), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_1005(1), ZN => gl_rom_n_1058);
  gl_rom_g35622 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_256(0), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_259(0), ZN => gl_rom_n_1057);
  gl_rom_g35623 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_1004(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_1003(1), ZN => gl_rom_n_1056);
  gl_rom_g35624 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_948(0), B1 => FE_OFN11_gl_rom_n_19, B2 => gl_rom_rom_946(0), ZN => gl_rom_n_1055);
  gl_rom_g35625 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_1000(1), B1 => FE_OFN19_gl_rom_n_16, B2 => gl_rom_rom_1006(1), ZN => gl_rom_n_1054);
  gl_rom_g35626 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_753(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_757(0), ZN => gl_rom_n_1053);
  gl_rom_g35627 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_985(1), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_989(1), ZN => gl_rom_n_1052);
  gl_rom_g35628 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_988(1), B1 => FE_OFN21_gl_rom_n_16, B2 => gl_rom_rom_990(1), ZN => gl_rom_n_1051);
  gl_rom_g35629 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_838(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_839(0), ZN => gl_rom_n_1050);
  gl_rom_g35630 : AOI22D0BWP7T port map(A1 => FE_OFN21_gl_rom_n_16, A2 => gl_rom_rom_374(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_375(0), ZN => gl_rom_n_1049);
  gl_rom_g35631 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_986(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_987(1), ZN => gl_rom_n_1048);
  gl_rom_g35632 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_984(1), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_991(1), ZN => gl_rom_n_1047);
  gl_rom_g35633 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_836(0), B1 => FE_OFN11_gl_rom_n_19, B2 => gl_rom_rom_834(0), ZN => gl_rom_n_1046);
  gl_rom_g35634 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_372(0), B1 => FE_OFN13_gl_rom_n_19, B2 => gl_rom_rom_370(0), ZN => gl_rom_n_1045);
  gl_rom_g35635 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_994(1), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_999(1), ZN => gl_rom_n_1044);
  gl_rom_g35636 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_996(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_998(1), ZN => gl_rom_n_1043);
  gl_rom_g35637 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_369(0), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_373(0), ZN => gl_rom_n_1042);
  gl_rom_g35638 : AOI22D0BWP7T port map(A1 => FE_OFN15_gl_rom_n_22, A2 => gl_rom_rom_997(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_995(1), ZN => gl_rom_n_1041);
  gl_rom_g35639 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_368(0), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_371(0), ZN => gl_rom_n_1040);
  gl_rom_g35640 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_992(1), B1 => FE_OFN25_gl_rom_n_21, B2 => gl_rom_rom_993(1), ZN => gl_rom_n_1039);
  gl_rom_g35641 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_833(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_837(0), ZN => gl_rom_n_1038);
  gl_rom_g35642 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_1010(1), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_1015(1), ZN => gl_rom_n_1037);
  gl_rom_g35643 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_752(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_755(0), ZN => gl_rom_n_1036);
  gl_rom_g35644 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_1012(1), B1 => FE_OFN21_gl_rom_n_16, B2 => gl_rom_rom_1014(1), ZN => gl_rom_n_1035);
  gl_rom_g35645 : AOI22D0BWP7T port map(A1 => FE_OFN21_gl_rom_n_16, A2 => gl_rom_rom_342(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_343(0), ZN => gl_rom_n_1034);
  gl_rom_g35646 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_832(0), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_835(0), ZN => gl_rom_n_1033);
  gl_rom_g35647 : AOI22D0BWP7T port map(A1 => FE_OFN15_gl_rom_n_22, A2 => gl_rom_rom_1013(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_1011(1), ZN => gl_rom_n_1032);
  gl_rom_g35648 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_1008(1), B1 => FE_OFN25_gl_rom_n_21, B2 => gl_rom_rom_1009(1), ZN => gl_rom_n_1031);
  gl_rom_g35649 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_340(0), B1 => FE_OFN13_gl_rom_n_19, B2 => gl_rom_rom_338(0), ZN => gl_rom_n_1030);
  gl_rom_g35650 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_978(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_983(1), ZN => gl_rom_n_1029);
  gl_rom_g35651 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_980(1), B1 => FE_OFN21_gl_rom_n_16, B2 => gl_rom_rom_982(1), ZN => gl_rom_n_1028);
  gl_rom_g35652 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_337(0), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_341(0), ZN => gl_rom_n_1027);
  gl_rom_g35653 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_977(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_981(0), ZN => gl_rom_n_1026);
  gl_rom_g35654 : AOI22D0BWP7T port map(A1 => FE_OFN15_gl_rom_n_22, A2 => gl_rom_rom_981(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_979(1), ZN => gl_rom_n_1025);
  gl_rom_g35655 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_336(0), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_339(0), ZN => gl_rom_n_1024);
  gl_rom_g35656 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_976(1), B1 => FE_OFN26_gl_rom_n_21, B2 => gl_rom_rom_977(1), ZN => gl_rom_n_1023);
  gl_rom_g35657 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_945(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_949(0), ZN => gl_rom_n_1022);
  gl_rom_g35658 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_969(1), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_973(1), ZN => gl_rom_n_1021);
  gl_rom_g35659 : AOI22D0BWP7T port map(A1 => FE_OFN17_gl_rom_n_16, A2 => gl_rom_rom_726(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_727(0), ZN => gl_rom_n_1020);
  gl_rom_g35660 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_972(1), B1 => FE_OFN21_gl_rom_n_16, B2 => gl_rom_rom_974(1), ZN => gl_rom_n_1019);
  gl_rom_g35661 : AOI22D0BWP7T port map(A1 => FE_OFN21_gl_rom_n_16, A2 => gl_rom_rom_350(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_351(0), ZN => gl_rom_n_1018);
  gl_rom_g35662 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_970(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_971(1), ZN => gl_rom_n_1017);
  gl_rom_g35663 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_968(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_975(1), ZN => gl_rom_n_1016);
  gl_rom_g35664 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_348(0), B1 => FE_OFN13_gl_rom_n_19, B2 => gl_rom_rom_346(0), ZN => gl_rom_n_1015);
  gl_rom_g35665 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_638(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_639(0), ZN => gl_rom_n_1014);
  gl_rom_g35666 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_962(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_967(1), ZN => gl_rom_n_1013);
  gl_rom_g35667 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_345(0), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_349(0), ZN => gl_rom_n_1012);
  gl_rom_g35668 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_964(1), B1 => FE_OFN21_gl_rom_n_16, B2 => gl_rom_rom_966(1), ZN => gl_rom_n_1011);
  gl_rom_g35669 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_724(0), B1 => FE_OFN11_gl_rom_n_19, B2 => gl_rom_rom_722(0), ZN => gl_rom_n_1010);
  gl_rom_g35670 : AOI22D0BWP7T port map(A1 => FE_OFN15_gl_rom_n_22, A2 => gl_rom_rom_965(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_963(1), ZN => gl_rom_n_1009);
  gl_rom_g35671 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_960(1), B1 => FE_OFN26_gl_rom_n_21, B2 => gl_rom_rom_961(1), ZN => gl_rom_n_1008);
  gl_rom_g35672 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_344(0), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_347(0), ZN => gl_rom_n_1007);
  gl_rom_g35673 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_953(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_959(1), ZN => gl_rom_n_1006);
  gl_rom_g35674 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_636(0), B1 => FE_OFN11_gl_rom_n_19, B2 => gl_rom_rom_634(0), ZN => gl_rom_n_1005);
  gl_rom_g35675 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_944(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_947(0), ZN => gl_rom_n_1004);
  gl_rom_g35676 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_954(1), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_957(1), ZN => gl_rom_n_1003);
  gl_rom_g35677 : AOI22D0BWP7T port map(A1 => FE_OFN21_gl_rom_n_16, A2 => gl_rom_rom_358(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_359(0), ZN => gl_rom_n_1002);
  gl_rom_g35678 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_956(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_958(1), ZN => gl_rom_n_1001);
  gl_rom_g35679 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_633(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_637(0), ZN => gl_rom_n_1000);
  gl_rom_g35680 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_356(0), B1 => FE_OFN12_gl_rom_n_19, B2 => gl_rom_rom_354(0), ZN => gl_rom_n_999);
  gl_rom_g35681 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_952(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_955(1), ZN => gl_rom_n_998);
  gl_rom_g35682 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_632(0), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_635(0), ZN => gl_rom_n_997);
  gl_rom_g35683 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_937(1), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_941(1), ZN => gl_rom_n_996);
  gl_rom_g35684 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_353(0), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_357(0), ZN => gl_rom_n_995);
  gl_rom_g35685 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_940(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_942(1), ZN => gl_rom_n_994);
  gl_rom_g35686 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_938(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_943(1), ZN => gl_rom_n_993);
  gl_rom_g35687 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_936(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_939(1), ZN => gl_rom_n_992);
  gl_rom_g35688 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_946(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_951(1), ZN => gl_rom_n_991);
  gl_rom_g35689 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_352(0), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_355(0), ZN => gl_rom_n_990);
  gl_rom_g35690 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_945(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_949(1), ZN => gl_rom_n_989);
  gl_rom_g35691 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_721(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_725(0), ZN => gl_rom_n_988);
  gl_rom_g35692 : AOI22D0BWP7T port map(A1 => FE_OFN21_gl_rom_n_16, A2 => gl_rom_rom_382(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_383(0), ZN => gl_rom_n_987);
  gl_rom_g35693 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_948(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_947(1), ZN => gl_rom_n_986);
  gl_rom_g35694 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_622(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_623(0), ZN => gl_rom_n_985);
  gl_rom_g35695 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_944(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_950(1), ZN => gl_rom_n_984);
  gl_rom_g35696 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_380(0), B1 => FE_OFN12_gl_rom_n_19, B2 => gl_rom_rom_378(0), ZN => gl_rom_n_983);
  gl_rom_g35697 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_720(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_723(0), ZN => gl_rom_n_982);
  gl_rom_g35698 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_914(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_919(1), ZN => gl_rom_n_981);
  gl_rom_g35699 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_913(1), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_917(1), ZN => gl_rom_n_980);
  gl_rom_g35700 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_377(0), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_381(0), ZN => gl_rom_n_979);
  gl_rom_g35701 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_916(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_915(1), ZN => gl_rom_n_978);
  gl_rom_g35702 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_376(0), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_379(0), ZN => gl_rom_n_977);
  gl_rom_g35703 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_912(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_918(1), ZN => gl_rom_n_976);
  gl_rom_g35704 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_620(0), B1 => FE_OFN11_gl_rom_n_19, B2 => gl_rom_rom_618(0), ZN => gl_rom_n_975);
  gl_rom_g35705 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_922(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_927(1), ZN => gl_rom_n_974);
  gl_rom_g35706 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_924(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_926(1), ZN => gl_rom_n_973);
  gl_rom_g35707 : AOI22D0BWP7T port map(A1 => FE_OFN21_gl_rom_n_16, A2 => gl_rom_rom_366(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_367(0), ZN => gl_rom_n_972);
  gl_rom_g35708 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_617(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_621(0), ZN => gl_rom_n_971);
  gl_rom_g35709 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_925(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_923(1), ZN => gl_rom_n_970);
  gl_rom_g35710 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_364(0), B1 => FE_OFN13_gl_rom_n_19, B2 => gl_rom_rom_362(0), ZN => gl_rom_n_969);
  gl_rom_g35711 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_920(1), B1 => FE_OFN26_gl_rom_n_21, B2 => gl_rom_rom_921(1), ZN => gl_rom_n_968);
  gl_rom_g35712 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_929(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_933(1), ZN => gl_rom_n_967);
  gl_rom_g35713 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_976(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_979(0), ZN => gl_rom_n_966);
  gl_rom_g35714 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_616(0), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_619(0), ZN => gl_rom_n_965);
  gl_rom_g35715 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_361(0), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_365(0), ZN => gl_rom_n_964);
  gl_rom_g35716 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_932(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_934(1), ZN => gl_rom_n_963);
  gl_rom_g35717 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_360(0), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_363(0), ZN => gl_rom_n_962);
  gl_rom_g35718 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_930(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_931(1), ZN => gl_rom_n_961);
  gl_rom_g35719 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_928(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_935(1), ZN => gl_rom_n_960);
  gl_rom_g35720 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_905(1), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_909(1), ZN => gl_rom_n_959);
  gl_rom_g35721 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_908(1), B1 => FE_OFN19_gl_rom_n_16, B2 => gl_rom_rom_910(1), ZN => gl_rom_n_958);
  gl_rom_g35722 : AOI22D0BWP7T port map(A1 => FE_OFN21_gl_rom_n_16, A2 => gl_rom_rom_334(0), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_335(0), ZN => gl_rom_n_957);
  gl_rom_g35723 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_729(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_733(0), ZN => gl_rom_n_956);
  gl_rom_g35724 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_906(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_911(1), ZN => gl_rom_n_955);
  gl_rom_g35725 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_904(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_907(1), ZN => gl_rom_n_954);
  gl_rom_g35726 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_332(0), B1 => FE_OFN12_gl_rom_n_19, B2 => gl_rom_rom_330(0), ZN => gl_rom_n_953);
  gl_rom_g35727 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_914(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_919(0), ZN => gl_rom_n_952);
  gl_rom_g35728 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_898(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_903(1), ZN => gl_rom_n_951);
  gl_rom_g35729 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_630(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_631(0), ZN => gl_rom_n_950);
  gl_rom_g35730 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_329(0), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_333(0), ZN => gl_rom_n_949);
  gl_rom_g35731 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_897(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_901(1), ZN => gl_rom_n_948);
  gl_rom_g35732 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_628(0), B1 => FE_OFN13_gl_rom_n_19, B2 => gl_rom_rom_626(0), ZN => gl_rom_n_947);
  gl_rom_g35733 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_328(0), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_331(0), ZN => gl_rom_n_946);
  gl_rom_g35734 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_900(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_899(1), ZN => gl_rom_n_945);
  gl_rom_g35735 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_896(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_902(1), ZN => gl_rom_n_944);
  gl_rom_g35736 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_732(0), B1 => FE_OFN17_gl_rom_n_16, B2 => gl_rom_rom_734(0), ZN => gl_rom_n_943);
  gl_rom_g35737 : AOI22D0BWP7T port map(A1 => FE_OFN21_gl_rom_n_16, A2 => gl_rom_rom_694(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_695(1), ZN => gl_rom_n_942);
  gl_rom_g35738 : AOI22D0BWP7T port map(A1 => FE_OFN21_gl_rom_n_16, A2 => gl_rom_rom_326(0), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_327(0), ZN => gl_rom_n_941);
  gl_rom_g35739 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_692(1), B1 => FE_OFN13_gl_rom_n_19, B2 => gl_rom_rom_690(1), ZN => gl_rom_n_940);
  gl_rom_g35740 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_625(0), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_629(0), ZN => gl_rom_n_939);
  gl_rom_g35741 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_689(1), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_693(1), ZN => gl_rom_n_938);
  gl_rom_g35742 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_688(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_691(1), ZN => gl_rom_n_937);
  gl_rom_g35743 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_324(0), B1 => FE_OFN12_gl_rom_n_19, B2 => gl_rom_rom_322(0), ZN => gl_rom_n_936);
  gl_rom_g35744 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_321(0), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_325(0), ZN => gl_rom_n_935);
  gl_rom_g35745 : AOI22D0BWP7T port map(A1 => FE_OFN21_gl_rom_n_16, A2 => gl_rom_rom_662(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_663(1), ZN => gl_rom_n_934);
  gl_rom_g35746 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_624(0), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_627(0), ZN => gl_rom_n_933);
  gl_rom_g35747 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_660(1), B1 => FE_OFN13_gl_rom_n_19, B2 => gl_rom_rom_658(1), ZN => gl_rom_n_932);
  gl_rom_g35748 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_320(0), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_323(0), ZN => gl_rom_n_931);
  gl_rom_g35749 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_657(1), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_661(1), ZN => gl_rom_n_930);
  gl_rom_g35750 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_656(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_659(1), ZN => gl_rom_n_929);
  gl_rom_g35751 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_730(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_731(0), ZN => gl_rom_n_928);
  gl_rom_g35752 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_665(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_671(1), ZN => gl_rom_n_927);
  gl_rom_g35753 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_666(1), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_669(1), ZN => gl_rom_n_926);
  gl_rom_g35754 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_913(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_917(0), ZN => gl_rom_n_925);
  gl_rom_g35755 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_122(0), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_127(0), ZN => gl_rom_n_924);
  gl_rom_g35756 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_668(1), B1 => FE_OFN21_gl_rom_n_16, B2 => gl_rom_rom_670(1), ZN => gl_rom_n_923);
  gl_rom_g35757 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_664(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_667(1), ZN => gl_rom_n_922);
  gl_rom_g35758 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_593(0), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_597(0), ZN => gl_rom_n_921);
  gl_rom_g35759 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_124(0), B1 => FE_OFN21_gl_rom_n_16, B2 => gl_rom_rom_126(0), ZN => gl_rom_n_920);
  gl_rom_g35760 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_674(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_679(1), ZN => gl_rom_n_919);
  gl_rom_g35761 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_728(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_735(0), ZN => gl_rom_n_918);
  gl_rom_g35762 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_673(1), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_677(1), ZN => gl_rom_n_917);
  gl_rom_g35763 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_596(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_598(0), ZN => gl_rom_n_916);
  gl_rom_g35764 : AOI22D0BWP7T port map(A1 => FE_OFN16_gl_rom_n_22, A2 => gl_rom_rom_125(0), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_123(0), ZN => gl_rom_n_915);
  gl_rom_g35765 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_120(0), B1 => FE_OFN26_gl_rom_n_21, B2 => gl_rom_rom_121(0), ZN => gl_rom_n_914);
  gl_rom_g35766 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_676(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_675(1), ZN => gl_rom_n_913);
  gl_rom_g35767 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_672(1), B1 => FE_OFN21_gl_rom_n_16, B2 => gl_rom_rom_678(1), ZN => gl_rom_n_912);
  gl_rom_g35768 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_697(1), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_701(1), ZN => gl_rom_n_911);
  gl_rom_g35769 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_1002(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_1007(0), ZN => gl_rom_n_910);
  gl_rom_g35770 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_594(0), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_595(0), ZN => gl_rom_n_909);
  gl_rom_g35771 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_700(1), B1 => FE_OFN21_gl_rom_n_16, B2 => gl_rom_rom_702(1), ZN => gl_rom_n_908);
  gl_rom_g35772 : AOI22D0BWP7T port map(A1 => FE_OFN21_gl_rom_n_16, A2 => gl_rom_rom_110(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_111(0), ZN => gl_rom_n_907);
  gl_rom_g35773 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_108(0), B1 => FE_OFN13_gl_rom_n_19, B2 => gl_rom_rom_106(0), ZN => gl_rom_n_906);
  gl_rom_g35774 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_698(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_699(1), ZN => gl_rom_n_905);
  gl_rom_g35775 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_696(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_703(1), ZN => gl_rom_n_904);
  gl_rom_g35776 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_681(1), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_685(1), ZN => gl_rom_n_903);
  gl_rom_g35777 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_592(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_599(0), ZN => gl_rom_n_902);
  gl_rom_g35778 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_105(0), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_109(0), ZN => gl_rom_n_901);
  gl_rom_g35779 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_684(1), B1 => FE_OFN21_gl_rom_n_16, B2 => gl_rom_rom_686(1), ZN => gl_rom_n_900);
  gl_rom_g35780 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_916(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_915(0), ZN => gl_rom_n_899);
  gl_rom_g35781 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_682(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_683(1), ZN => gl_rom_n_898);
  gl_rom_g35782 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_104(0), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_107(0), ZN => gl_rom_n_897);
  gl_rom_g35783 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_680(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_687(1), ZN => gl_rom_n_896);
  gl_rom_g35784 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_737(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_743(0), ZN => gl_rom_n_895);
  gl_rom_g35785 : AOI22D0BWP7T port map(A1 => FE_OFN21_gl_rom_n_16, A2 => gl_rom_rom_654(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_655(1), ZN => gl_rom_n_894);
  gl_rom_g35786 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_652(1), B1 => FE_OFN13_gl_rom_n_19, B2 => gl_rom_rom_650(1), ZN => gl_rom_n_893);
  gl_rom_g35787 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_89(0), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_93(0), ZN => gl_rom_n_892);
  gl_rom_g35788 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_649(1), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_653(1), ZN => gl_rom_n_891);
  gl_rom_g35789 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_92(0), B1 => FE_OFN21_gl_rom_n_16, B2 => gl_rom_rom_94(0), ZN => gl_rom_n_890);
  gl_rom_g35790 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_648(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_651(1), ZN => gl_rom_n_889);
  gl_rom_g35791 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_606(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_607(0), ZN => gl_rom_n_888);
  gl_rom_g35792 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_604(0), B1 => FE_OFN11_gl_rom_n_19, B2 => gl_rom_rom_602(0), ZN => gl_rom_n_887);
  gl_rom_g35793 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_642(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_647(1), ZN => gl_rom_n_886);
  gl_rom_g35794 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_90(0), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_91(0), ZN => gl_rom_n_885);
  gl_rom_g35795 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_644(1), B1 => FE_OFN21_gl_rom_n_16, B2 => gl_rom_rom_646(1), ZN => gl_rom_n_884);
  gl_rom_g35796 : AOI22D0BWP7T port map(A1 => FE_OFN15_gl_rom_n_22, A2 => gl_rom_rom_645(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_643(1), ZN => gl_rom_n_883);
  gl_rom_g35797 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_640(1), B1 => FE_OFN26_gl_rom_n_21, B2 => gl_rom_rom_641(1), ZN => gl_rom_n_882);
  gl_rom_g35798 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_562(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_567(1), ZN => gl_rom_n_881);
  gl_rom_g35799 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_88(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_95(0), ZN => gl_rom_n_880);
  gl_rom_g35800 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_738(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_741(0), ZN => gl_rom_n_879);
  gl_rom_g35801 : AOI22D0BWP7T port map(A1 => FE_OFN21_gl_rom_n_16, A2 => gl_rom_rom_102(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_103(0), ZN => gl_rom_n_878);
  gl_rom_g35802 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_564(1), B1 => FE_OFN21_gl_rom_n_16, B2 => gl_rom_rom_566(1), ZN => gl_rom_n_877);
  gl_rom_g35803 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_601(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_605(0), ZN => gl_rom_n_876);
  gl_rom_g35804 : AOI22D0BWP7T port map(A1 => FE_OFN15_gl_rom_n_22, A2 => gl_rom_rom_565(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_563(1), ZN => gl_rom_n_875);
  gl_rom_g35805 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_100(0), B1 => FE_OFN12_gl_rom_n_19, B2 => gl_rom_rom_98(0), ZN => gl_rom_n_874);
  gl_rom_g35806 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_560(1), B1 => FE_OFN26_gl_rom_n_21, B2 => gl_rom_rom_561(1), ZN => gl_rom_n_873);
  gl_rom_g35807 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_985(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_989(0), ZN => gl_rom_n_872);
  gl_rom_g35808 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_97(0), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_101(0), ZN => gl_rom_n_871);
  gl_rom_g35809 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_530(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_535(1), ZN => gl_rom_n_870);
  gl_rom_g35810 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_600(0), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_603(0), ZN => gl_rom_n_869);
  gl_rom_g35811 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_532(1), B1 => FE_OFN21_gl_rom_n_16, B2 => gl_rom_rom_534(1), ZN => gl_rom_n_868);
  gl_rom_g35812 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_912(0), B1 => FE_OFN17_gl_rom_n_16, B2 => gl_rom_rom_918(0), ZN => gl_rom_n_867);
  gl_rom_g35813 : AOI22D0BWP7T port map(A1 => FE_OFN15_gl_rom_n_22, A2 => gl_rom_rom_533(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_531(1), ZN => gl_rom_n_866);
  gl_rom_g35814 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_96(0), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_99(0), ZN => gl_rom_n_865);
  gl_rom_g35815 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_528(1), B1 => FE_OFN26_gl_rom_n_21, B2 => gl_rom_rom_529(1), ZN => gl_rom_n_864);
  gl_rom_g35816 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_740(0), B1 => FE_OFN17_gl_rom_n_16, B2 => gl_rom_rom_742(0), ZN => gl_rom_n_863);
  gl_rom_g35817 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_537(1), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_541(1), ZN => gl_rom_n_862);
  gl_rom_g35818 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_1004(0), B1 => FE_OFN17_gl_rom_n_16, B2 => gl_rom_rom_1006(0), ZN => gl_rom_n_861);
  gl_rom_g35819 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_736(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_739(0), ZN => gl_rom_n_860);
  gl_rom_g35820 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_540(1), B1 => FE_OFN21_gl_rom_n_16, B2 => gl_rom_rom_542(1), ZN => gl_rom_n_859);
  gl_rom_g35821 : AOI22D0BWP7T port map(A1 => FE_OFN21_gl_rom_n_16, A2 => gl_rom_rom_118(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_119(0), ZN => gl_rom_n_858);
  gl_rom_g35822 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_614(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_615(0), ZN => gl_rom_n_857);
  gl_rom_g35823 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_538(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_539(1), ZN => gl_rom_n_856);
  gl_rom_g35824 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_116(0), B1 => FE_OFN12_gl_rom_n_19, B2 => gl_rom_rom_114(0), ZN => gl_rom_n_855);
  gl_rom_g35825 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_536(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_543(1), ZN => gl_rom_n_854);
  gl_rom_g35826 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_546(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_551(1), ZN => gl_rom_n_853);
  gl_rom_g35827 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_113(0), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_117(0), ZN => gl_rom_n_852);
  gl_rom_g35828 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_548(1), B1 => FE_OFN21_gl_rom_n_16, B2 => gl_rom_rom_550(1), ZN => gl_rom_n_851);
  gl_rom_g35829 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_612(0), B1 => FE_OFN11_gl_rom_n_19, B2 => gl_rom_rom_610(0), ZN => gl_rom_n_850);
  gl_rom_g35830 : AOI22D0BWP7T port map(A1 => FE_OFN15_gl_rom_n_22, A2 => gl_rom_rom_549(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_547(1), ZN => gl_rom_n_849);
  gl_rom_g35831 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_544(1), B1 => FE_OFN26_gl_rom_n_21, B2 => gl_rom_rom_545(1), ZN => gl_rom_n_848);
  gl_rom_g35832 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_112(0), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_115(0), ZN => gl_rom_n_847);
  gl_rom_g35833 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_569(1), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_573(1), ZN => gl_rom_n_846);
  gl_rom_g35834 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_609(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_613(0), ZN => gl_rom_n_845);
  gl_rom_g35835 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_16, A2 => gl_rom_rom_86(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_87(0), ZN => gl_rom_n_844);
  gl_rom_g35836 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_572(1), B1 => FE_OFN19_gl_rom_n_16, B2 => gl_rom_rom_574(1), ZN => gl_rom_n_843);
  gl_rom_g35837 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_84(0), B1 => FE_OFN12_gl_rom_n_19, B2 => gl_rom_rom_82(0), ZN => gl_rom_n_842);
  gl_rom_g35838 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_570(1), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_575(1), ZN => gl_rom_n_841);
  gl_rom_g35839 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_568(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_571(1), ZN => gl_rom_n_840);
  gl_rom_g35840 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_16, A2 => gl_rom_rom_558(1), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_559(1), ZN => gl_rom_n_839);
  gl_rom_g35841 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_608(0), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_611(0), ZN => gl_rom_n_838);
  gl_rom_g35842 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_81(0), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_85(0), ZN => gl_rom_n_837);
  gl_rom_g35843 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_556(1), B1 => FE_OFN13_gl_rom_n_19, B2 => gl_rom_rom_554(1), ZN => gl_rom_n_836);
  gl_rom_g35844 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_80(0), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_83(0), ZN => gl_rom_n_835);
  gl_rom_g35845 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_553(1), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_557(1), ZN => gl_rom_n_834);
  gl_rom_g35846 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_552(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_555(1), ZN => gl_rom_n_833);
  gl_rom_g35847 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_522(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_527(1), ZN => gl_rom_n_832);
  gl_rom_g35848 : AOI22D0BWP7T port map(A1 => FE_OFN17_gl_rom_n_16, A2 => gl_rom_rom_718(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_719(0), ZN => gl_rom_n_831);
  gl_rom_g35849 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_524(1), B1 => FE_OFN21_gl_rom_n_16, B2 => gl_rom_rom_526(1), ZN => gl_rom_n_830);
  gl_rom_g35850 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_16, A2 => gl_rom_rom_78(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_79(0), ZN => gl_rom_n_829);
  gl_rom_g35851 : AOI22D0BWP7T port map(A1 => FE_OFN15_gl_rom_n_22, A2 => gl_rom_rom_525(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_523(1), ZN => gl_rom_n_828);
  gl_rom_g35852 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_590(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_591(0), ZN => gl_rom_n_827);
  gl_rom_g35853 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_520(1), B1 => FE_OFN26_gl_rom_n_21, B2 => gl_rom_rom_521(1), ZN => gl_rom_n_826);
  gl_rom_g35854 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_76(0), B1 => FE_OFN12_gl_rom_n_19, B2 => gl_rom_rom_74(0), ZN => gl_rom_n_825);
  gl_rom_g35855 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_926(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_927(0), ZN => gl_rom_n_824);
  gl_rom_g35856 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_514(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_519(1), ZN => gl_rom_n_823);
  gl_rom_g35857 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_73(0), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_77(0), ZN => gl_rom_n_822);
  gl_rom_g35858 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_516(1), B1 => FE_OFN21_gl_rom_n_16, B2 => gl_rom_rom_518(1), ZN => gl_rom_n_821);
  gl_rom_g35859 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_72(0), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_75(0), ZN => gl_rom_n_820);
  gl_rom_g35860 : AOI22D0BWP7T port map(A1 => FE_OFN15_gl_rom_n_22, A2 => gl_rom_rom_517(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_515(1), ZN => gl_rom_n_819);
  gl_rom_g35861 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_512(1), B1 => FE_OFN26_gl_rom_n_21, B2 => gl_rom_rom_513(1), ZN => gl_rom_n_818);
  gl_rom_g35862 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_588(0), B1 => FE_OFN13_gl_rom_n_19, B2 => gl_rom_rom_586(0), ZN => gl_rom_n_817);
  gl_rom_g35863 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_988(0), B1 => FE_OFN17_gl_rom_n_16, B2 => gl_rom_rom_990(0), ZN => gl_rom_n_816);
  gl_rom_g35864 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_16, A2 => gl_rom_rom_70(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_71(0), ZN => gl_rom_n_815);
  gl_rom_g35865 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_585(0), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_589(0), ZN => gl_rom_n_814);
  gl_rom_g35866 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_506(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_511(1), ZN => gl_rom_n_813);
  gl_rom_g35867 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_505(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_509(1), ZN => gl_rom_n_812);
  gl_rom_g35868 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_716(0), B1 => FE_OFN11_gl_rom_n_19, B2 => gl_rom_rom_714(0), ZN => gl_rom_n_811);
  gl_rom_g35869 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_68(0), B1 => FE_OFN12_gl_rom_n_19, B2 => gl_rom_rom_66(0), ZN => gl_rom_n_810);
  gl_rom_g35870 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_508(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_507(1), ZN => gl_rom_n_809);
  gl_rom_g35871 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_504(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_510(1), ZN => gl_rom_n_808);
  gl_rom_g35872 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_65(0), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_69(0), ZN => gl_rom_n_807);
  gl_rom_g35873 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_1016(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_1019(1), ZN => gl_rom_n_806);
  gl_rom_g35874 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_64(0), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_67(0), ZN => gl_rom_n_805);
  gl_rom_g35875 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_490(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_495(1), ZN => gl_rom_n_804);
  gl_rom_g35876 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_489(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_493(1), ZN => gl_rom_n_803);
  gl_rom_g35877 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_713(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_717(0), ZN => gl_rom_n_802);
  gl_rom_g35878 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_492(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_491(1), ZN => gl_rom_n_801);
  gl_rom_g35879 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_488(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_494(1), ZN => gl_rom_n_800);
  gl_rom_g35880 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_474(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_479(1), ZN => gl_rom_n_799);
  gl_rom_g35881 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_924(0), B1 => FE_OFN11_gl_rom_n_19, B2 => gl_rom_rom_922(0), ZN => gl_rom_n_798);
  gl_rom_g35882 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_582(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_583(0), ZN => gl_rom_n_797);
  gl_rom_g35883 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_476(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_478(1), ZN => gl_rom_n_796);
  gl_rom_g35884 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_16, A2 => gl_rom_rom_510(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_511(0), ZN => gl_rom_n_795);
  gl_rom_g35885 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_477(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_475(1), ZN => gl_rom_n_794);
  gl_rom_g35886 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_472(1), B1 => FE_OFN26_gl_rom_n_21, B2 => gl_rom_rom_473(1), ZN => gl_rom_n_793);
  gl_rom_g35887 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_508(0), B1 => FE_OFN13_gl_rom_n_19, B2 => gl_rom_rom_506(0), ZN => gl_rom_n_792);
  gl_rom_g35888 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_580(0), B1 => FE_OFN13_gl_rom_n_19, B2 => gl_rom_rom_578(0), ZN => gl_rom_n_791);
  gl_rom_g35889 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_481(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_485(1), ZN => gl_rom_n_790);
  gl_rom_g35890 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_484(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_486(1), ZN => gl_rom_n_789);
  gl_rom_g35891 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_505(0), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_509(0), ZN => gl_rom_n_788);
  gl_rom_g35892 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_482(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_483(1), ZN => gl_rom_n_787);
  gl_rom_g35893 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_480(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_487(1), ZN => gl_rom_n_786);
  gl_rom_g35894 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_504(0), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_507(0), ZN => gl_rom_n_785);
  gl_rom_g35895 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_497(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_501(1), ZN => gl_rom_n_784);
  gl_rom_g35896 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_712(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_715(0), ZN => gl_rom_n_783);
  gl_rom_g35897 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_577(0), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_581(0), ZN => gl_rom_n_782);
  gl_rom_g35898 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_489(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_495(0), ZN => gl_rom_n_781);
  gl_rom_g35899 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_500(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_502(1), ZN => gl_rom_n_780);
  gl_rom_g35900 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_498(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_499(1), ZN => gl_rom_n_779);
  gl_rom_g35901 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_576(0), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_579(0), ZN => gl_rom_n_778);
  gl_rom_g35902 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_496(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_503(1), ZN => gl_rom_n_777);
  gl_rom_g35903 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_490(0), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_493(0), ZN => gl_rom_n_776);
  gl_rom_g35904 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_465(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_469(1), ZN => gl_rom_n_775);
  gl_rom_g35905 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_492(0), B1 => FE_OFN19_gl_rom_n_16, B2 => gl_rom_rom_494(0), ZN => gl_rom_n_774);
  gl_rom_g35906 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_468(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_470(1), ZN => gl_rom_n_773);
  gl_rom_g35907 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_466(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_471(1), ZN => gl_rom_n_772);
  gl_rom_g35908 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_1020(0), B1 => FE_OFN17_gl_rom_n_16, B2 => gl_rom_rom_1022(0), ZN => gl_rom_n_771);
  gl_rom_g35909 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_710(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_711(0), ZN => gl_rom_n_770);
  gl_rom_g35910 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_488(0), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_491(0), ZN => gl_rom_n_769);
  gl_rom_g35911 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_464(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_467(1), ZN => gl_rom_n_768);
  gl_rom_g35912 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_921(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_925(0), ZN => gl_rom_n_767);
  gl_rom_g35913 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_457(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_461(1), ZN => gl_rom_n_766);
  gl_rom_g35914 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_460(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_462(1), ZN => gl_rom_n_765);
  gl_rom_g35915 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_474(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_479(0), ZN => gl_rom_n_764);
  gl_rom_g35916 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_458(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_459(1), ZN => gl_rom_n_763);
  gl_rom_g35917 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_456(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_463(1), ZN => gl_rom_n_762);
  gl_rom_g35918 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_476(0), B1 => FE_OFN19_gl_rom_n_16, B2 => gl_rom_rom_478(0), ZN => gl_rom_n_761);
  gl_rom_g35919 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_708(0), B1 => FE_OFN11_gl_rom_n_19, B2 => gl_rom_rom_706(0), ZN => gl_rom_n_760);
  gl_rom_g35920 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_697(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_701(0), ZN => gl_rom_n_759);
  gl_rom_g35921 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_450(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_455(1), ZN => gl_rom_n_758);
  gl_rom_g35922 : AOI22D0BWP7T port map(A1 => FE_OFN15_gl_rom_n_22, A2 => gl_rom_rom_477(0), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_475(0), ZN => gl_rom_n_757);
  gl_rom_g35923 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_452(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_454(1), ZN => gl_rom_n_756);
  gl_rom_g35924 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_986(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_987(0), ZN => gl_rom_n_755);
  gl_rom_g35925 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_453(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_451(1), ZN => gl_rom_n_754);
  gl_rom_g35926 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_472(0), B1 => FE_OFN26_gl_rom_n_21, B2 => gl_rom_rom_473(0), ZN => gl_rom_n_753);
  gl_rom_g35927 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_448(1), B1 => gl_rom_n_21, B2 => gl_rom_rom_449(1), ZN => gl_rom_n_752);
  gl_rom_g35928 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_700(0), B1 => FE_OFN17_gl_rom_n_16, B2 => gl_rom_rom_702(0), ZN => gl_rom_n_751);
  gl_rom_g35929 : AOI22D0BWP7T port map(A1 => FE_OFN14_gl_rom_n_22, A2 => gl_rom_rom_1005(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_1003(0), ZN => gl_rom_n_750);
  gl_rom_g35930 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_441(1), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_445(1), ZN => gl_rom_n_749);
  gl_rom_g35931 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_481(0), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_485(0), ZN => gl_rom_n_748);
  gl_rom_g35932 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_444(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_446(1), ZN => gl_rom_n_747);
  gl_rom_g35933 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_484(0), B1 => FE_OFN19_gl_rom_n_16, B2 => gl_rom_rom_486(0), ZN => gl_rom_n_746);
  gl_rom_g35934 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_442(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_443(1), ZN => gl_rom_n_745);
  gl_rom_g35935 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_440(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_447(1), ZN => gl_rom_n_744);
  gl_rom_g35936 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_698(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_699(0), ZN => gl_rom_n_743);
  gl_rom_g35937 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_920(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_923(0), ZN => gl_rom_n_742);
  gl_rom_g35938 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_705(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_709(0), ZN => gl_rom_n_741);
  gl_rom_g35939 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_16, A2 => gl_rom_rom_430(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_431(1), ZN => gl_rom_n_740);
  gl_rom_g35940 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_482(0), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_483(0), ZN => gl_rom_n_739);
  gl_rom_g35941 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_428(1), B1 => FE_OFN12_gl_rom_n_19, B2 => gl_rom_rom_426(1), ZN => gl_rom_n_738);
  gl_rom_g35942 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_425(1), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_429(1), ZN => gl_rom_n_737);
  gl_rom_g35943 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_424(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_427(1), ZN => gl_rom_n_736);
  gl_rom_g35944 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_480(0), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_487(0), ZN => gl_rom_n_735);
  gl_rom_g35945 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_704(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_707(0), ZN => gl_rom_n_734);
  gl_rom_g35946 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_409(1), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_413(1), ZN => gl_rom_n_733);
  gl_rom_g35947 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_412(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_414(1), ZN => gl_rom_n_732);
  gl_rom_g35948 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_696(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_703(0), ZN => gl_rom_n_731);
  gl_rom_g35949 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_16, A2 => gl_rom_rom_502(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_503(0), ZN => gl_rom_n_730);
  gl_rom_g35950 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_410(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_411(1), ZN => gl_rom_n_729);
  gl_rom_g35951 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_408(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_415(1), ZN => gl_rom_n_728);
  gl_rom_g35952 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_500(0), B1 => FE_OFN12_gl_rom_n_19, B2 => gl_rom_rom_498(0), ZN => gl_rom_n_727);
  gl_rom_g35953 : AOI22D0BWP7T port map(A1 => FE_OFN17_gl_rom_n_16, A2 => gl_rom_rom_686(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_687(0), ZN => gl_rom_n_726);
  gl_rom_g35954 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_417(1), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_421(1), ZN => gl_rom_n_725);
  gl_rom_g35955 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_497(0), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_501(0), ZN => gl_rom_n_724);
  gl_rom_g35956 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_420(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_422(1), ZN => gl_rom_n_723);
  gl_rom_g35957 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_684(0), B1 => gl_rom_n_19, B2 => gl_rom_rom_682(0), ZN => gl_rom_n_722);
  gl_rom_g35958 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_418(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_423(1), ZN => gl_rom_n_721);
  gl_rom_g35959 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_416(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_419(1), ZN => gl_rom_n_720);
  gl_rom_g35960 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_496(0), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_499(0), ZN => gl_rom_n_719);
  gl_rom_g35961 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_433(1), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_437(1), ZN => gl_rom_n_718);
  gl_rom_g35962 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_436(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_438(1), ZN => gl_rom_n_717);
  gl_rom_g35963 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_465(0), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_469(0), ZN => gl_rom_n_716);
  gl_rom_g35964 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_434(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_435(1), ZN => gl_rom_n_715);
  gl_rom_g35965 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_468(0), B1 => FE_OFN19_gl_rom_n_16, B2 => gl_rom_rom_470(0), ZN => gl_rom_n_714);
  gl_rom_g35966 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_432(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_439(1), ZN => gl_rom_n_713);
  gl_rom_g35967 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_681(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_685(0), ZN => gl_rom_n_712);
  gl_rom_g35968 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_16, A2 => gl_rom_rom_406(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_407(1), ZN => gl_rom_n_711);
  gl_rom_g35969 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_466(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_471(0), ZN => gl_rom_n_710);
  gl_rom_g35970 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_404(1), B1 => FE_OFN12_gl_rom_n_19, B2 => gl_rom_rom_402(1), ZN => gl_rom_n_709);
  gl_rom_g35971 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_680(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_683(0), ZN => gl_rom_n_708);
  gl_rom_g35972 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_401(1), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_405(1), ZN => gl_rom_n_707);
  gl_rom_g35973 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_984(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_991(0), ZN => gl_rom_n_706);
  gl_rom_g35974 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_464(0), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_467(0), ZN => gl_rom_n_705);
  gl_rom_g35975 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_400(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_403(1), ZN => gl_rom_n_704);
  gl_rom_g35976 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_929(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_935(0), ZN => gl_rom_n_703);
  gl_rom_g35977 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_16, A2 => gl_rom_rom_398(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_399(1), ZN => gl_rom_n_702);
  gl_rom_g35978 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_396(1), B1 => FE_OFN12_gl_rom_n_19, B2 => gl_rom_rom_394(1), ZN => gl_rom_n_701);
  gl_rom_g35979 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_457(0), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_461(0), ZN => gl_rom_n_700);
  gl_rom_g35980 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_393(1), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_397(1), ZN => gl_rom_n_699);
  gl_rom_g35981 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_930(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_933(0), ZN => gl_rom_n_698);
  gl_rom_g35982 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_460(0), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_462(0), ZN => gl_rom_n_697);
  gl_rom_g35983 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_392(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_395(1), ZN => gl_rom_n_696);
  gl_rom_g35984 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_689(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_693(0), ZN => gl_rom_n_695);
  gl_rom_g35985 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_385(1), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_389(1), ZN => gl_rom_n_694);
  gl_rom_g35986 : AOI22D0BWP7T port map(A1 => FE_OFN17_gl_rom_n_16, A2 => gl_rom_rom_830(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_831(0), ZN => gl_rom_n_693);
  gl_rom_g35987 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_388(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_390(1), ZN => gl_rom_n_692);
  gl_rom_g35988 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_458(0), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_463(0), ZN => gl_rom_n_691);
  gl_rom_g35989 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_386(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_391(1), ZN => gl_rom_n_690);
  gl_rom_g35990 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_692(0), B1 => FE_OFN17_gl_rom_n_16, B2 => gl_rom_rom_694(0), ZN => gl_rom_n_689);
  gl_rom_g35991 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_456(0), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_459(0), ZN => gl_rom_n_688);
  gl_rom_g35992 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_384(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_387(1), ZN => gl_rom_n_687);
  gl_rom_g35993 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_449(0), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_455(0), ZN => gl_rom_n_686);
  gl_rom_g35994 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_378(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_383(1), ZN => gl_rom_n_685);
  gl_rom_g35995 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_380(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_382(1), ZN => gl_rom_n_684);
  gl_rom_g35996 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_690(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_691(0), ZN => gl_rom_n_683);
  gl_rom_g35997 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_450(0), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_453(0), ZN => gl_rom_n_682);
  gl_rom_g35998 : AOI22D0BWP7T port map(A1 => FE_OFN16_gl_rom_n_22, A2 => gl_rom_rom_381(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_379(1), ZN => gl_rom_n_681);
  gl_rom_g35999 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_376(1), B1 => FE_OFN27_gl_rom_n_21, B2 => gl_rom_rom_377(1), ZN => gl_rom_n_680);
  gl_rom_g36000 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_828(0), B1 => gl_rom_n_19, B2 => gl_rom_rom_826(0), ZN => gl_rom_n_679);
  gl_rom_g36001 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_452(0), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_454(0), ZN => gl_rom_n_678);
  gl_rom_g36002 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_362(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_367(1), ZN => gl_rom_n_677);
  gl_rom_g36003 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_364(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_366(1), ZN => gl_rom_n_676);
  gl_rom_g36004 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_448(0), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_451(0), ZN => gl_rom_n_675);
  gl_rom_g36005 : AOI22D0BWP7T port map(A1 => FE_OFN16_gl_rom_n_22, A2 => gl_rom_rom_365(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_363(1), ZN => gl_rom_n_674);
  gl_rom_g36006 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_360(1), B1 => FE_OFN27_gl_rom_n_21, B2 => gl_rom_rom_361(1), ZN => gl_rom_n_673);
  gl_rom_g36007 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_688(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_695(0), ZN => gl_rom_n_672);
  gl_rom_g36008 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_370(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_375(1), ZN => gl_rom_n_671);
  gl_rom_g36009 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_369(1), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_373(1), ZN => gl_rom_n_670);
  gl_rom_g36010 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_825(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_829(0), ZN => gl_rom_n_669);
  gl_rom_g36011 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_441(0), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_445(0), ZN => gl_rom_n_668);
  gl_rom_g36012 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_372(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_371(1), ZN => gl_rom_n_667);
  gl_rom_g36013 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_368(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_374(1), ZN => gl_rom_n_666);
  gl_rom_g36014 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_657(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_661(0), ZN => gl_rom_n_665);
  gl_rom_g36015 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_444(0), B1 => FE_OFN19_gl_rom_n_16, B2 => gl_rom_rom_446(0), ZN => gl_rom_n_664);
  gl_rom_g36016 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_660(0), B1 => FE_OFN17_gl_rom_n_16, B2 => gl_rom_rom_662(0), ZN => gl_rom_n_663);
  gl_rom_g36017 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_337(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_343(1), ZN => gl_rom_n_662);
  gl_rom_g36018 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_338(1), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_341(1), ZN => gl_rom_n_661);
  gl_rom_g36019 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_442(0), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_443(0), ZN => gl_rom_n_660);
  gl_rom_g36020 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_340(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_342(1), ZN => gl_rom_n_659);
  gl_rom_g36021 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_336(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_339(1), ZN => gl_rom_n_658);
  gl_rom_g36022 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_440(0), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_447(0), ZN => gl_rom_n_657);
  gl_rom_g36023 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_346(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_351(1), ZN => gl_rom_n_656);
  gl_rom_g36024 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_658(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_659(0), ZN => gl_rom_n_655);
  gl_rom_g36025 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_348(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_350(1), ZN => gl_rom_n_654);
  gl_rom_g36026 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_425(0), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_431(0), ZN => gl_rom_n_653);
  gl_rom_g36027 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_824(0), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_827(0), ZN => gl_rom_n_652);
  gl_rom_g36028 : AOI22D0BWP7T port map(A1 => FE_OFN15_gl_rom_n_22, A2 => gl_rom_rom_349(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_347(1), ZN => gl_rom_n_651);
  gl_rom_g36029 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_426(0), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_429(0), ZN => gl_rom_n_650);
  gl_rom_g36030 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_344(1), B1 => FE_OFN27_gl_rom_n_21, B2 => gl_rom_rom_345(1), ZN => gl_rom_n_649);
  gl_rom_g36031 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_656(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_663(0), ZN => gl_rom_n_648);
  gl_rom_g36032 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_354(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_359(1), ZN => gl_rom_n_647);
  gl_rom_g36033 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_353(1), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_357(1), ZN => gl_rom_n_646);
  gl_rom_g36034 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_428(0), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_430(0), ZN => gl_rom_n_645);
  gl_rom_g36035 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_356(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_355(1), ZN => gl_rom_n_644);
  gl_rom_g36036 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_424(0), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_427(0), ZN => gl_rom_n_643);
  gl_rom_g36037 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_352(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_358(1), ZN => gl_rom_n_642);
  gl_rom_g36038 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_1000(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_1001(0), ZN => gl_rom_n_641);
  gl_rom_g36039 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_330(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_335(1), ZN => gl_rom_n_640);
  gl_rom_g36040 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_932(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_934(0), ZN => gl_rom_n_639);
  gl_rom_g36041 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_332(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_334(1), ZN => gl_rom_n_638);
  gl_rom_g36042 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_433(0), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_437(0), ZN => gl_rom_n_637);
  gl_rom_g36043 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_928(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_931(0), ZN => gl_rom_n_636);
  gl_rom_g36044 : AOI22D0BWP7T port map(A1 => FE_OFN15_gl_rom_n_22, A2 => gl_rom_rom_333(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_331(1), ZN => gl_rom_n_635);
  gl_rom_g36045 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_328(1), B1 => FE_OFN26_gl_rom_n_21, B2 => gl_rom_rom_329(1), ZN => gl_rom_n_634);
  gl_rom_g36046 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_436(0), B1 => FE_OFN19_gl_rom_n_16, B2 => gl_rom_rom_438(0), ZN => gl_rom_n_633);
  gl_rom_g36047 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_665(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_669(0), ZN => gl_rom_n_632);
  gl_rom_g36048 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_322(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_327(1), ZN => gl_rom_n_631);
  gl_rom_g36049 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_434(0), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_435(0), ZN => gl_rom_n_630);
  gl_rom_g36050 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_321(1), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_325(1), ZN => gl_rom_n_629);
  gl_rom_g36051 : AOI22D0BWP7T port map(A1 => FE_OFN17_gl_rom_n_16, A2 => gl_rom_rom_814(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_815(0), ZN => gl_rom_n_628);
  gl_rom_g36052 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_432(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_439(0), ZN => gl_rom_n_627);
  gl_rom_g36053 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_324(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_323(1), ZN => gl_rom_n_626);
  gl_rom_g36054 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_320(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_326(1), ZN => gl_rom_n_625);
  gl_rom_g36055 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_668(0), B1 => FE_OFN17_gl_rom_n_16, B2 => gl_rom_rom_670(0), ZN => gl_rom_n_624);
  gl_rom_g36056 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_812(0), B1 => gl_rom_n_19, B2 => gl_rom_rom_810(0), ZN => gl_rom_n_623);
  gl_rom_g36057 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_122(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_127(1), ZN => gl_rom_n_622);
  gl_rom_g36058 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_402(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_407(0), ZN => gl_rom_n_621);
  gl_rom_g36059 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_124(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_126(1), ZN => gl_rom_n_620);
  gl_rom_g36060 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_666(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_667(0), ZN => gl_rom_n_619);
  gl_rom_g36061 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_404(0), B1 => FE_OFN19_gl_rom_n_16, B2 => gl_rom_rom_406(0), ZN => gl_rom_n_618);
  gl_rom_g36062 : AOI22D0BWP7T port map(A1 => FE_OFN15_gl_rom_n_22, A2 => gl_rom_rom_125(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_123(1), ZN => gl_rom_n_617);
  gl_rom_g36063 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_664(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_671(0), ZN => gl_rom_n_616);
  gl_rom_g36064 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_120(1), B1 => FE_OFN26_gl_rom_n_21, B2 => gl_rom_rom_121(1), ZN => gl_rom_n_615);
  gl_rom_g36065 : AOI22D0BWP7T port map(A1 => FE_OFN15_gl_rom_n_22, A2 => gl_rom_rom_405(0), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_403(0), ZN => gl_rom_n_614);
  gl_rom_g36066 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_106(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_111(1), ZN => gl_rom_n_613);
  gl_rom_g36067 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_108(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_110(1), ZN => gl_rom_n_612);
  gl_rom_g36068 : AOI22D0BWP7T port map(A1 => FE_OFN15_gl_rom_n_22, A2 => gl_rom_rom_109(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_107(1), ZN => gl_rom_n_611);
  gl_rom_g36069 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_104(1), B1 => FE_OFN27_gl_rom_n_21, B2 => gl_rom_rom_105(1), ZN => gl_rom_n_610);
  gl_rom_g36070 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_400(0), B1 => FE_OFN26_gl_rom_n_21, B2 => gl_rom_rom_401(0), ZN => gl_rom_n_609);
  gl_rom_g36071 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_809(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_813(0), ZN => gl_rom_n_608);
  gl_rom_g36072 : AOI22D0BWP7T port map(A1 => FE_OFN21_gl_rom_n_16, A2 => gl_rom_rom_118(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_119(1), ZN => gl_rom_n_607);
  gl_rom_g36073 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_116(1), B1 => FE_OFN12_gl_rom_n_19, B2 => gl_rom_rom_114(1), ZN => gl_rom_n_606);
  gl_rom_g36074 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_16, A2 => gl_rom_rom_414(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_415(0), ZN => gl_rom_n_605);
  gl_rom_g36075 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_993(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_999(0), ZN => gl_rom_n_604);
  gl_rom_g36076 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_113(1), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_117(1), ZN => gl_rom_n_603);
  gl_rom_g36077 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_112(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_115(1), ZN => gl_rom_n_602);
  gl_rom_g36078 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_412(0), B1 => FE_OFN12_gl_rom_n_19, B2 => gl_rom_rom_410(0), ZN => gl_rom_n_601);
  gl_rom_g36079 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_673(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_677(0), ZN => gl_rom_n_600);
  gl_rom_g36080 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_81(1), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_85(1), ZN => gl_rom_n_599);
  gl_rom_g36081 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_409(0), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_413(0), ZN => gl_rom_n_598);
  gl_rom_g36082 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_84(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_86(1), ZN => gl_rom_n_597);
  gl_rom_g36083 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_676(0), B1 => FE_OFN17_gl_rom_n_16, B2 => gl_rom_rom_678(0), ZN => gl_rom_n_596);
  gl_rom_g36084 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_82(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_83(1), ZN => gl_rom_n_595);
  gl_rom_g36085 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_80(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_87(1), ZN => gl_rom_n_594);
  gl_rom_g36086 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_408(0), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_411(0), ZN => gl_rom_n_593);
  gl_rom_g36087 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_90(1), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_95(1), ZN => gl_rom_n_592);
  gl_rom_g36088 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_417(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_423(0), ZN => gl_rom_n_591);
  gl_rom_g36089 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_92(1), B1 => FE_OFN21_gl_rom_n_16, B2 => gl_rom_rom_94(1), ZN => gl_rom_n_590);
  gl_rom_g36090 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_808(0), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_811(0), ZN => gl_rom_n_589);
  gl_rom_g36091 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_674(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_675(0), ZN => gl_rom_n_588);
  gl_rom_g36092 : AOI22D0BWP7T port map(A1 => FE_OFN15_gl_rom_n_22, A2 => gl_rom_rom_93(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_91(1), ZN => gl_rom_n_587);
  gl_rom_g36093 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_88(1), B1 => FE_OFN26_gl_rom_n_21, B2 => gl_rom_rom_89(1), ZN => gl_rom_n_586);
  gl_rom_g36094 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_418(0), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_421(0), ZN => gl_rom_n_585);
  gl_rom_g36095 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_420(0), B1 => FE_OFN19_gl_rom_n_16, B2 => gl_rom_rom_422(0), ZN => gl_rom_n_584);
  gl_rom_g36096 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_97(1), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_101(1), ZN => gl_rom_n_583);
  gl_rom_g36097 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_100(1), B1 => FE_OFN21_gl_rom_n_16, B2 => gl_rom_rom_102(1), ZN => gl_rom_n_582);
  gl_rom_g36098 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_672(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_679(0), ZN => gl_rom_n_581);
  gl_rom_g36099 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_98(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_99(1), ZN => gl_rom_n_580);
  gl_rom_g36100 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_416(0), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_419(0), ZN => gl_rom_n_579);
  gl_rom_g36101 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_96(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_103(1), ZN => gl_rom_n_578);
  gl_rom_g36102 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_994(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_997(0), ZN => gl_rom_n_577);
  gl_rom_g36103 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_74(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_79(1), ZN => gl_rom_n_576);
  gl_rom_g36104 : AOI22D0BWP7T port map(A1 => FE_OFN17_gl_rom_n_16, A2 => gl_rom_rom_958(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_959(0), ZN => gl_rom_n_575);
  gl_rom_g36105 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_393(0), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_399(0), ZN => gl_rom_n_574);
  gl_rom_g36106 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_76(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_78(1), ZN => gl_rom_n_573);
  gl_rom_g36107 : AOI22D0BWP7T port map(A1 => FE_OFN15_gl_rom_n_22, A2 => gl_rom_rom_77(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_75(1), ZN => gl_rom_n_572);
  gl_rom_g36108 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_649(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_653(0), ZN => gl_rom_n_571);
  gl_rom_g36109 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_394(0), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_397(0), ZN => gl_rom_n_570);
  gl_rom_g36110 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_72(1), B1 => FE_OFN26_gl_rom_n_21, B2 => gl_rom_rom_73(1), ZN => gl_rom_n_569);
  gl_rom_g36111 : AOI22D0BWP7T port map(A1 => FE_OFN17_gl_rom_n_16, A2 => gl_rom_rom_822(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_823(0), ZN => gl_rom_n_568);
  gl_rom_g36112 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_65(1), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_69(1), ZN => gl_rom_n_567);
  gl_rom_g36113 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_396(0), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_398(0), ZN => gl_rom_n_566);
  gl_rom_g36114 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_68(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_70(1), ZN => gl_rom_n_565);
  gl_rom_g36115 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_392(0), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_395(0), ZN => gl_rom_n_564);
  gl_rom_g36116 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_66(1), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_67(1), ZN => gl_rom_n_563);
  gl_rom_g36117 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_64(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_71(1), ZN => gl_rom_n_562);
  gl_rom_g36118 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_652(0), B1 => FE_OFN17_gl_rom_n_16, B2 => gl_rom_rom_654(0), ZN => gl_rom_n_561);
  gl_rom_g36119 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_16, A2 => gl_rom_rom_390(0), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_391(0), ZN => gl_rom_n_560);
  gl_rom_g36120 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_218(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_223(1), ZN => gl_rom_n_559);
  gl_rom_g36121 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_820(0), B1 => FE_OFN11_gl_rom_n_19, B2 => gl_rom_rom_818(0), ZN => gl_rom_n_558);
  gl_rom_g36122 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_220(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_222(1), ZN => gl_rom_n_557);
  gl_rom_g36123 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_388(0), B1 => FE_OFN12_gl_rom_n_19, B2 => gl_rom_rom_386(0), ZN => gl_rom_n_556);
  gl_rom_g36124 : AOI22D0BWP7T port map(A1 => FE_OFN16_gl_rom_n_22, A2 => gl_rom_rom_221(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_219(1), ZN => gl_rom_n_555);
  gl_rom_g36125 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_650(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_651(0), ZN => gl_rom_n_554);
  gl_rom_g36126 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_216(1), B1 => FE_OFN27_gl_rom_n_21, B2 => gl_rom_rom_217(1), ZN => gl_rom_n_553);
  gl_rom_g36127 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_385(0), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_389(0), ZN => gl_rom_n_552);
  gl_rom_g36128 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_648(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_655(0), ZN => gl_rom_n_551);
  gl_rom_g36129 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_756(1), B1 => FE_OFN19_gl_rom_n_16, B2 => gl_rom_rom_758(1), ZN => gl_rom_n_550);
  gl_rom_g36130 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_226(1), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_229(1), ZN => gl_rom_n_549);
  gl_rom_g36131 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_384(0), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_387(0), ZN => gl_rom_n_548);
  gl_rom_g36132 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_228(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_230(1), ZN => gl_rom_n_547);
  gl_rom_g36133 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_224(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_227(1), ZN => gl_rom_n_546);
  gl_rom_g36134 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_956(0), B1 => FE_OFN11_gl_rom_n_19, B2 => gl_rom_rom_954(0), ZN => gl_rom_n_545);
  gl_rom_g36135 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_242(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_247(1), ZN => gl_rom_n_544);
  gl_rom_g36136 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_244(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_246(1), ZN => gl_rom_n_543);
  gl_rom_g36137 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_817(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_821(0), ZN => gl_rom_n_542);
  gl_rom_g36138 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_185(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_189(0), ZN => gl_rom_n_541);
  gl_rom_g36139 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_641(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_645(0), ZN => gl_rom_n_540);
  gl_rom_g36140 : AOI22D0BWP7T port map(A1 => FE_OFN16_gl_rom_n_22, A2 => gl_rom_rom_245(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_243(1), ZN => gl_rom_n_539);
  gl_rom_g36141 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_188(0), B1 => FE_OFN17_gl_rom_n_16, B2 => gl_rom_rom_190(0), ZN => gl_rom_n_538);
  gl_rom_g36142 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_240(1), B1 => FE_OFN27_gl_rom_n_21, B2 => gl_rom_rom_241(1), ZN => gl_rom_n_537);
  gl_rom_g36143 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_210(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_215(1), ZN => gl_rom_n_536);
  gl_rom_g36144 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_186(0), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_187(0), ZN => gl_rom_n_535);
  gl_rom_g36145 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_212(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_214(1), ZN => gl_rom_n_534);
  gl_rom_g36146 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_644(0), B1 => FE_OFN17_gl_rom_n_16, B2 => gl_rom_rom_646(0), ZN => gl_rom_n_533);
  gl_rom_g36147 : AOI22D0BWP7T port map(A1 => FE_OFN16_gl_rom_n_22, A2 => gl_rom_rom_213(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_211(1), ZN => gl_rom_n_532);
  gl_rom_g36148 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_184(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_191(0), ZN => gl_rom_n_531);
  gl_rom_g36149 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_208(1), B1 => FE_OFN27_gl_rom_n_21, B2 => gl_rom_rom_209(1), ZN => gl_rom_n_530);
  gl_rom_g36150 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_816(0), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_819(0), ZN => gl_rom_n_529);
  gl_rom_g36151 : AOI22D0BWP7T port map(A1 => FE_OFN21_gl_rom_n_16, A2 => gl_rom_rom_254(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_255(1), ZN => gl_rom_n_528);
  gl_rom_g36152 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_642(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_643(0), ZN => gl_rom_n_527);
  gl_rom_g36153 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_252(1), B1 => FE_OFN12_gl_rom_n_19, B2 => gl_rom_rom_250(1), ZN => gl_rom_n_526);
  gl_rom_g36154 : AOI22D0BWP7T port map(A1 => FE_OFN17_gl_rom_n_16, A2 => gl_rom_rom_174(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_175(0), ZN => gl_rom_n_525);
  gl_rom_g36155 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_172(0), B1 => gl_rom_n_19, B2 => gl_rom_rom_170(0), ZN => gl_rom_n_524);
  gl_rom_g36156 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_249(1), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_253(1), ZN => gl_rom_n_523);
  gl_rom_g36157 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_248(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_251(1), ZN => gl_rom_n_522);
  gl_rom_g36158 : AOI22D0BWP7T port map(A1 => FE_OFN21_gl_rom_n_16, A2 => gl_rom_rom_238(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_239(1), ZN => gl_rom_n_521);
  gl_rom_g36159 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_640(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_647(0), ZN => gl_rom_n_520);
  gl_rom_g36160 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_169(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_173(0), ZN => gl_rom_n_519);
  gl_rom_g36161 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_236(1), B1 => FE_OFN12_gl_rom_n_19, B2 => gl_rom_rom_234(1), ZN => gl_rom_n_518);
  gl_rom_g36162 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_168(0), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_171(0), ZN => gl_rom_n_517);
  gl_rom_g36163 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_233(1), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_237(1), ZN => gl_rom_n_516);
  gl_rom_g36164 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_232(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_235(1), ZN => gl_rom_n_515);
  gl_rom_g36165 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_953(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_957(0), ZN => gl_rom_n_514);
  gl_rom_g36166 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_201(1), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_205(1), ZN => gl_rom_n_513);
  gl_rom_g36167 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_204(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_206(1), ZN => gl_rom_n_512);
  gl_rom_g36168 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_178(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_183(0), ZN => gl_rom_n_511);
  gl_rom_g36169 : AOI22D0BWP7T port map(A1 => FE_OFN17_gl_rom_n_16, A2 => gl_rom_rom_790(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_791(0), ZN => gl_rom_n_510);
  gl_rom_g36170 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_202(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_203(1), ZN => gl_rom_n_509);
  gl_rom_g36171 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_200(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_207(1), ZN => gl_rom_n_508);
  gl_rom_g36172 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_177(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_181(0), ZN => gl_rom_n_507);
  gl_rom_g36173 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_16, A2 => gl_rom_rom_198(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_199(1), ZN => gl_rom_n_506);
  gl_rom_g36174 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_569(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_573(0), ZN => gl_rom_n_505);
  gl_rom_g36175 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_180(0), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_179(0), ZN => gl_rom_n_504);
  gl_rom_g36176 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_196(1), B1 => FE_OFN12_gl_rom_n_19, B2 => gl_rom_rom_194(1), ZN => gl_rom_n_503);
  gl_rom_g36177 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_572(0), B1 => FE_OFN17_gl_rom_n_16, B2 => gl_rom_rom_574(0), ZN => gl_rom_n_502);
  gl_rom_g36178 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_176(0), B1 => FE_OFN17_gl_rom_n_16, B2 => gl_rom_rom_182(0), ZN => gl_rom_n_501);
  gl_rom_g36179 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_193(1), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_197(1), ZN => gl_rom_n_500);
  gl_rom_g36180 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_192(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_195(1), ZN => gl_rom_n_499);
  gl_rom_g36181 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_788(0), B1 => FE_OFN11_gl_rom_n_19, B2 => gl_rom_rom_786(0), ZN => gl_rom_n_498);
  gl_rom_g36182 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_306(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_311(1), ZN => gl_rom_n_497);
  gl_rom_g36183 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_146(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_151(0), ZN => gl_rom_n_496);
  gl_rom_g36184 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_308(1), B1 => FE_OFN21_gl_rom_n_16, B2 => gl_rom_rom_310(1), ZN => gl_rom_n_495);
  gl_rom_g36185 : AOI22D0BWP7T port map(A1 => FE_OFN16_gl_rom_n_22, A2 => gl_rom_rom_309(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_307(1), ZN => gl_rom_n_494);
  gl_rom_g36186 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_570(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_571(0), ZN => gl_rom_n_493);
  gl_rom_g36187 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_148(0), B1 => FE_OFN17_gl_rom_n_16, B2 => gl_rom_rom_150(0), ZN => gl_rom_n_492);
  gl_rom_g36188 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_304(1), B1 => FE_OFN27_gl_rom_n_21, B2 => gl_rom_rom_305(1), ZN => gl_rom_n_491);
  gl_rom_g36189 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_952(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_955(0), ZN => gl_rom_n_490);
  gl_rom_g36190 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_274(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_279(1), ZN => gl_rom_n_489);
  gl_rom_g36191 : AOI22D0BWP7T port map(A1 => FE_OFN14_gl_rom_n_22, A2 => gl_rom_rom_149(0), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_147(0), ZN => gl_rom_n_488);
  gl_rom_g36192 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_568(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_575(0), ZN => gl_rom_n_487);
  gl_rom_g36193 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_276(1), B1 => FE_OFN21_gl_rom_n_16, B2 => gl_rom_rom_278(1), ZN => gl_rom_n_486);
  gl_rom_g36194 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_144(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_145(0), ZN => gl_rom_n_485);
  gl_rom_g36195 : AOI22D0BWP7T port map(A1 => FE_OFN16_gl_rom_n_22, A2 => gl_rom_rom_277(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_275(1), ZN => gl_rom_n_484);
  gl_rom_g36196 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_272(1), B1 => FE_OFN27_gl_rom_n_21, B2 => gl_rom_rom_273(1), ZN => gl_rom_n_483);
  gl_rom_g36197 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_996(0), B1 => FE_OFN17_gl_rom_n_16, B2 => gl_rom_rom_998(0), ZN => gl_rom_n_482);
  gl_rom_g36198 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_282(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_287(1), ZN => gl_rom_n_481);
  gl_rom_g36199 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_785(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_789(0), ZN => gl_rom_n_480);
  gl_rom_g36200 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_284(1), B1 => FE_OFN21_gl_rom_n_16, B2 => gl_rom_rom_286(1), ZN => gl_rom_n_479);
  gl_rom_g36201 : AOI22D0BWP7T port map(A1 => FE_OFN17_gl_rom_n_16, A2 => gl_rom_rom_158(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_159(0), ZN => gl_rom_n_478);
  gl_rom_g36202 : AOI22D0BWP7T port map(A1 => FE_OFN16_gl_rom_n_22, A2 => gl_rom_rom_285(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_283(1), ZN => gl_rom_n_477);
  gl_rom_g36203 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_784(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_787(0), ZN => gl_rom_n_476);
  gl_rom_g36204 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_156(0), B1 => FE_OFN11_gl_rom_n_19, B2 => gl_rom_rom_154(0), ZN => gl_rom_n_475);
  gl_rom_g36205 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_280(1), B1 => FE_OFN27_gl_rom_n_21, B2 => gl_rom_rom_281(1), ZN => gl_rom_n_474);
  gl_rom_g36206 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_553(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_557(0), ZN => gl_rom_n_473);
  gl_rom_g36207 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_290(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_295(1), ZN => gl_rom_n_472);
  gl_rom_g36208 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_556(0), B1 => FE_OFN17_gl_rom_n_16, B2 => gl_rom_rom_558(0), ZN => gl_rom_n_471);
  gl_rom_g36209 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_292(1), B1 => FE_OFN21_gl_rom_n_16, B2 => gl_rom_rom_294(1), ZN => gl_rom_n_470);
  gl_rom_g36210 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_153(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_157(0), ZN => gl_rom_n_469);
  gl_rom_g36211 : AOI22D0BWP7T port map(A1 => FE_OFN16_gl_rom_n_22, A2 => gl_rom_rom_293(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_291(1), ZN => gl_rom_n_468);
  gl_rom_g36212 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_152(0), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_155(0), ZN => gl_rom_n_467);
  gl_rom_g36213 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_288(1), B1 => FE_OFN27_gl_rom_n_21, B2 => gl_rom_rom_289(1), ZN => gl_rom_n_466);
  gl_rom_g36214 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_313(1), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_317(1), ZN => gl_rom_n_465);
  gl_rom_g36215 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_161(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_165(0), ZN => gl_rom_n_464);
  gl_rom_g36216 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_316(1), B1 => FE_OFN21_gl_rom_n_16, B2 => gl_rom_rom_318(1), ZN => gl_rom_n_463);
  gl_rom_g36217 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_554(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_555(0), ZN => gl_rom_n_462);
  gl_rom_g36218 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_314(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_315(1), ZN => gl_rom_n_461);
  gl_rom_g36219 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_164(0), B1 => FE_OFN17_gl_rom_n_16, B2 => gl_rom_rom_166(0), ZN => gl_rom_n_460);
  gl_rom_g36220 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_312(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_319(1), ZN => gl_rom_n_459);
  gl_rom_g36221 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_297(1), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_301(1), ZN => gl_rom_n_458);
  gl_rom_g36222 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_162(0), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_163(0), ZN => gl_rom_n_457);
  gl_rom_g36223 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_300(1), B1 => FE_OFN21_gl_rom_n_16, B2 => gl_rom_rom_302(1), ZN => gl_rom_n_456);
  gl_rom_g36224 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_992(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_995(0), ZN => gl_rom_n_455);
  gl_rom_g36225 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_552(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_559(0), ZN => gl_rom_n_454);
  gl_rom_g36226 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_298(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_299(1), ZN => gl_rom_n_453);
  gl_rom_g36227 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_160(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_167(0), ZN => gl_rom_n_452);
  gl_rom_g36228 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_296(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_303(1), ZN => gl_rom_n_451);
  gl_rom_g36229 : AOI22D0BWP7T port map(A1 => FE_OFN17_gl_rom_n_16, A2 => gl_rom_rom_942(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_943(0), ZN => gl_rom_n_450);
  gl_rom_g36230 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_265(1), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_269(1), ZN => gl_rom_n_449);
  gl_rom_g36231 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_137(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_141(0), ZN => gl_rom_n_448);
  gl_rom_g36232 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_268(1), B1 => FE_OFN21_gl_rom_n_16, B2 => gl_rom_rom_270(1), ZN => gl_rom_n_447);
  gl_rom_g36233 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_266(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_267(1), ZN => gl_rom_n_446);
  gl_rom_g36234 : AOI22D0BWP7T port map(A1 => FE_OFN17_gl_rom_n_16, A2 => gl_rom_rom_798(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_799(0), ZN => gl_rom_n_445);
  gl_rom_g36235 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_140(0), B1 => FE_OFN17_gl_rom_n_16, B2 => gl_rom_rom_142(0), ZN => gl_rom_n_444);
  gl_rom_g36236 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_264(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_271(1), ZN => gl_rom_n_443);
  gl_rom_g36237 : AOI22D0BWP7T port map(A1 => FE_OFN17_gl_rom_n_16, A2 => gl_rom_rom_566(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_567(0), ZN => gl_rom_n_442);
  gl_rom_g36238 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_258(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_263(1), ZN => gl_rom_n_441);
  gl_rom_g36239 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_138(0), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_139(0), ZN => gl_rom_n_440);
  gl_rom_g36240 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_260(1), B1 => FE_OFN21_gl_rom_n_16, B2 => gl_rom_rom_262(1), ZN => gl_rom_n_439);
  gl_rom_g36241 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_136(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_143(0), ZN => gl_rom_n_438);
  gl_rom_g36242 : AOI22D0BWP7T port map(A1 => FE_OFN16_gl_rom_n_22, A2 => gl_rom_rom_261(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_259(1), ZN => gl_rom_n_437);
  gl_rom_g36243 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_256(1), B1 => FE_OFN27_gl_rom_n_21, B2 => gl_rom_rom_257(1), ZN => gl_rom_n_436);
  gl_rom_g36244 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_564(0), B1 => gl_rom_n_19, B2 => gl_rom_rom_562(0), ZN => gl_rom_n_435);
  gl_rom_g36245 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_130(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_135(0), ZN => gl_rom_n_434);
  gl_rom_g36246 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_186(1), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_191(1), ZN => gl_rom_n_433);
  gl_rom_g36247 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_796(0), B1 => gl_rom_n_19, B2 => gl_rom_rom_794(0), ZN => gl_rom_n_432);
  gl_rom_g36248 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_188(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_190(1), ZN => gl_rom_n_431);
  gl_rom_g36249 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_129(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_133(0), ZN => gl_rom_n_430);
  gl_rom_g36250 : AOI22D0BWP7T port map(A1 => FE_OFN14_gl_rom_n_22, A2 => gl_rom_rom_189(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_187(1), ZN => gl_rom_n_429);
  gl_rom_g36251 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_561(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_565(0), ZN => gl_rom_n_428);
  gl_rom_g36252 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_184(1), B1 => FE_OFN25_gl_rom_n_21, B2 => gl_rom_rom_185(1), ZN => gl_rom_n_427);
  gl_rom_g36253 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_132(0), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_131(0), ZN => gl_rom_n_426);
  gl_rom_g36254 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_1009(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_1013(0), ZN => gl_rom_n_425);
  gl_rom_g36255 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_560(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_563(0), ZN => gl_rom_n_424);
  gl_rom_g36256 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_170(1), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_175(1), ZN => gl_rom_n_423);
  gl_rom_g36257 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_172(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_174(1), ZN => gl_rom_n_422);
  gl_rom_g36258 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_128(0), B1 => FE_OFN17_gl_rom_n_16, B2 => gl_rom_rom_134(0), ZN => gl_rom_n_421);
  gl_rom_g36259 : AOI22D0BWP7T port map(A1 => FE_OFN14_gl_rom_n_22, A2 => gl_rom_rom_173(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_171(1), ZN => gl_rom_n_420);
  gl_rom_g36260 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_940(0), B1 => FE_OFN11_gl_rom_n_19, B2 => gl_rom_rom_938(0), ZN => gl_rom_n_419);
  gl_rom_g36261 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_168(1), B1 => FE_OFN25_gl_rom_n_21, B2 => gl_rom_rom_169(1), ZN => gl_rom_n_418);
  gl_rom_g36262 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_177(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_181(1), ZN => gl_rom_n_417);
  gl_rom_g36263 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_793(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_797(0), ZN => gl_rom_n_416);
  gl_rom_g36264 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_180(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_182(1), ZN => gl_rom_n_415);
  gl_rom_g36265 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_62(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_63(0), ZN => gl_rom_n_414);
  gl_rom_g36266 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_178(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_179(1), ZN => gl_rom_n_413);
  gl_rom_g36267 : AOI22D0BWP7T port map(A1 => FE_OFN17_gl_rom_n_16, A2 => gl_rom_rom_534(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_535(0), ZN => gl_rom_n_412);
  gl_rom_g36268 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_176(1), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_183(1), ZN => gl_rom_n_411);
  gl_rom_g36269 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_60(0), B1 => FE_OFN11_gl_rom_n_19, B2 => gl_rom_rom_58(0), ZN => gl_rom_n_410);
  gl_rom_g36270 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_146(1), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_151(1), ZN => gl_rom_n_409);
  gl_rom_g36271 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_145(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_149(1), ZN => gl_rom_n_408);
  gl_rom_g36272 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_57(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_61(0), ZN => gl_rom_n_407);
  gl_rom_g36273 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_56(0), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_59(0), ZN => gl_rom_n_406);
  gl_rom_g36274 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_148(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_147(1), ZN => gl_rom_n_405);
  gl_rom_g36275 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_144(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_150(1), ZN => gl_rom_n_404);
  gl_rom_g36276 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_532(0), B1 => gl_rom_n_19, B2 => gl_rom_rom_530(0), ZN => gl_rom_n_403);
  gl_rom_g36277 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_154(1), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_159(1), ZN => gl_rom_n_402);
  gl_rom_g36278 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_792(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_795(0), ZN => gl_rom_n_401);
  gl_rom_g36279 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_46(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_47(0), ZN => gl_rom_n_400);
  gl_rom_g36280 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_156(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_158(1), ZN => gl_rom_n_399);
  gl_rom_g36281 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_529(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_533(0), ZN => gl_rom_n_398);
  gl_rom_g36282 : AOI22D0BWP7T port map(A1 => FE_OFN14_gl_rom_n_22, A2 => gl_rom_rom_157(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_155(1), ZN => gl_rom_n_397);
  gl_rom_g36283 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_44(0), B1 => FE_OFN11_gl_rom_n_19, B2 => gl_rom_rom_42(0), ZN => gl_rom_n_396);
  gl_rom_g36284 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_152(1), B1 => FE_OFN25_gl_rom_n_21, B2 => gl_rom_rom_153(1), ZN => gl_rom_n_395);
  gl_rom_g36285 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_162(1), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_167(1), ZN => gl_rom_n_394);
  gl_rom_g36286 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_528(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_531(0), ZN => gl_rom_n_393);
  gl_rom_g36287 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_41(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_45(0), ZN => gl_rom_n_392);
  gl_rom_g36288 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_164(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_166(1), ZN => gl_rom_n_391);
  gl_rom_g36289 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_40(0), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_43(0), ZN => gl_rom_n_390);
  gl_rom_g36290 : AOI22D0BWP7T port map(A1 => FE_OFN14_gl_rom_n_22, A2 => gl_rom_rom_165(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_163(1), ZN => gl_rom_n_389);
  gl_rom_g36291 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_160(1), B1 => FE_OFN25_gl_rom_n_21, B2 => gl_rom_rom_161(1), ZN => gl_rom_n_388);
  gl_rom_g36292 : AOI22D0BWP7T port map(A1 => FE_OFN14_gl_rom_n_22, A2 => gl_rom_rom_1021(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_1019(0), ZN => gl_rom_n_387);
  gl_rom_g36293 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_937(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_941(0), ZN => gl_rom_n_386);
  gl_rom_g36294 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_138(1), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_143(1), ZN => gl_rom_n_385);
  gl_rom_g36295 : AOI22D0BWP7T port map(A1 => FE_OFN17_gl_rom_n_16, A2 => gl_rom_rom_806(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_807(0), ZN => gl_rom_n_384);
  gl_rom_g36296 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_140(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_142(1), ZN => gl_rom_n_383);
  gl_rom_g36297 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_54(0), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_55(0), ZN => gl_rom_n_382);
  gl_rom_g36298 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_141(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_139(1), ZN => gl_rom_n_381);
  gl_rom_g36299 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_52(0), B1 => FE_OFN11_gl_rom_n_19, B2 => gl_rom_rom_50(0), ZN => gl_rom_n_380);
  gl_rom_g36300 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_136(1), B1 => FE_OFN25_gl_rom_n_21, B2 => gl_rom_rom_137(1), ZN => gl_rom_n_379);
  gl_rom_g36301 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_537(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_541(0), ZN => gl_rom_n_378);
  gl_rom_g36302 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_130(1), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_135(1), ZN => gl_rom_n_377);
  gl_rom_g36303 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_49(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_53(0), ZN => gl_rom_n_376);
  gl_rom_g36304 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_132(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_134(1), ZN => gl_rom_n_375);
  gl_rom_g36305 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_540(0), B1 => FE_OFN17_gl_rom_n_16, B2 => gl_rom_rom_542(0), ZN => gl_rom_n_374);
  gl_rom_g36306 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_48(0), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_51(0), ZN => gl_rom_n_373);
  gl_rom_g36307 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_133(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_131(1), ZN => gl_rom_n_372);
  gl_rom_g36308 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_128(1), B1 => FE_OFN25_gl_rom_n_21, B2 => gl_rom_rom_129(1), ZN => gl_rom_n_371);
  gl_rom_g36309 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_804(0), B1 => gl_rom_n_19, B2 => gl_rom_rom_802(0), ZN => gl_rom_n_370);
  gl_rom_g36310 : AOI22D0BWP7T port map(A1 => FE_OFN17_gl_rom_n_16, A2 => gl_rom_rom_62(1), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_63(1), ZN => gl_rom_n_369);
  gl_rom_g36311 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_17(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_21(0), ZN => gl_rom_n_368);
  gl_rom_g36312 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_60(1), B1 => FE_OFN11_gl_rom_n_19, B2 => gl_rom_rom_58(1), ZN => gl_rom_n_367);
  gl_rom_g36313 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_57(1), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_61(1), ZN => gl_rom_n_366);
  gl_rom_g36314 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_20(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_22(0), ZN => gl_rom_n_365);
  gl_rom_g36315 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_56(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_59(1), ZN => gl_rom_n_364);
  gl_rom_g36316 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_936(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_939(0), ZN => gl_rom_n_363);
  gl_rom_g36317 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_538(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_539(0), ZN => gl_rom_n_362);
  gl_rom_g36318 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_18(0), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_19(0), ZN => gl_rom_n_361);
  gl_rom_g36319 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_41(1), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_47(1), ZN => gl_rom_n_360);
  gl_rom_g36320 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_536(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_543(0), ZN => gl_rom_n_359);
  gl_rom_g36321 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_42(1), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_45(1), ZN => gl_rom_n_358);
  gl_rom_g36322 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_16(0), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_23(0), ZN => gl_rom_n_357);
  gl_rom_g36323 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_44(1), B1 => FE_OFN17_gl_rom_n_16, B2 => gl_rom_rom_46(1), ZN => gl_rom_n_356);
  gl_rom_g36324 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_40(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_43(1), ZN => gl_rom_n_355);
  gl_rom_g36325 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_25(1), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_29(1), ZN => gl_rom_n_354);
  gl_rom_g36326 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_801(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_805(0), ZN => gl_rom_n_353);
  gl_rom_g36327 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_30(0), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_31(0), ZN => gl_rom_n_352);
  gl_rom_g36328 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_28(1), B1 => FE_OFN17_gl_rom_n_16, B2 => gl_rom_rom_30(1), ZN => gl_rom_n_351);
  gl_rom_g36329 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_545(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_549(0), ZN => gl_rom_n_350);
  gl_rom_g36330 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_26(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_27(1), ZN => gl_rom_n_349);
  gl_rom_g36331 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_28(0), B1 => FE_OFN11_gl_rom_n_19, B2 => gl_rom_rom_26(0), ZN => gl_rom_n_348);
  gl_rom_g36332 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_24(1), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_31(1), ZN => gl_rom_n_347);
  gl_rom_g36333 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_33(1), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_37(1), ZN => gl_rom_n_346);
  gl_rom_g36334 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_969(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_975(0), ZN => gl_rom_n_345);
  gl_rom_g36335 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_36(1), B1 => FE_OFN17_gl_rom_n_16, B2 => gl_rom_rom_38(1), ZN => gl_rom_n_344);
  gl_rom_g36336 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_25(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_29(0), ZN => gl_rom_n_343);
  gl_rom_g36337 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_800(0), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_803(0), ZN => gl_rom_n_342);
  gl_rom_g36338 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_548(0), B1 => FE_OFN17_gl_rom_n_16, B2 => gl_rom_rom_550(0), ZN => gl_rom_n_341);
  gl_rom_g36339 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_34(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_35(1), ZN => gl_rom_n_340);
  gl_rom_g36340 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_24(0), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_27(0), ZN => gl_rom_n_339);
  gl_rom_g36341 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_32(1), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_39(1), ZN => gl_rom_n_338);
  gl_rom_g36342 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_50(1), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_55(1), ZN => gl_rom_n_337);
  gl_rom_g36343 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_33(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_37(0), ZN => gl_rom_n_336);
  gl_rom_g36344 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_52(1), B1 => FE_OFN17_gl_rom_n_16, B2 => gl_rom_rom_54(1), ZN => gl_rom_n_335);
  gl_rom_g36345 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_36(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_38(0), ZN => gl_rom_n_334);
  gl_rom_g36346 : AOI22D0BWP7T port map(A1 => FE_OFN14_gl_rom_n_22, A2 => gl_rom_rom_53(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_51(1), ZN => gl_rom_n_333);
  gl_rom_g36347 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_48(1), B1 => FE_OFN25_gl_rom_n_21, B2 => gl_rom_rom_49(1), ZN => gl_rom_n_332);
  gl_rom_g36348 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_546(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_547(0), ZN => gl_rom_n_331);
  gl_rom_g36349 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_18(1), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_23(1), ZN => gl_rom_n_330);
  gl_rom_g36350 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_544(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_551(0), ZN => gl_rom_n_329);
  gl_rom_g36351 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_34(0), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_35(0), ZN => gl_rom_n_328);
  gl_rom_g36352 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_20(1), B1 => FE_OFN17_gl_rom_n_16, B2 => gl_rom_rom_22(1), ZN => gl_rom_n_327);
  gl_rom_g36353 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_1012(0), B1 => FE_OFN17_gl_rom_n_16, B2 => gl_rom_rom_1014(0), ZN => gl_rom_n_326);
  gl_rom_g36354 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_32(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_39(0), ZN => gl_rom_n_325);
  gl_rom_g36355 : AOI22D0BWP7T port map(A1 => FE_OFN14_gl_rom_n_22, A2 => gl_rom_rom_21(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_19(1), ZN => gl_rom_n_324);
  gl_rom_g36356 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_16(1), B1 => gl_rom_n_21, B2 => gl_rom_rom_17(1), ZN => gl_rom_n_323);
  gl_rom_g36357 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_910(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_911(0), ZN => gl_rom_n_322);
  gl_rom_g36358 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_9(1), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_13(1), ZN => gl_rom_n_321);
  gl_rom_g36359 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_14(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_15(0), ZN => gl_rom_n_320);
  gl_rom_g36360 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_12(1), B1 => FE_OFN17_gl_rom_n_16, B2 => gl_rom_rom_14(1), ZN => gl_rom_n_319);
  gl_rom_g36361 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_10(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_11(1), ZN => gl_rom_n_318);
  gl_rom_g36362 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_777(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_781(0), ZN => gl_rom_n_317);
  gl_rom_g36363 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_12(0), B1 => FE_OFN11_gl_rom_n_19, B2 => gl_rom_rom_10(0), ZN => gl_rom_n_316);
  gl_rom_g36364 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_8(1), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_15(1), ZN => gl_rom_n_315);
  gl_rom_g36365 : AOI22D0BWP7T port map(A1 => FE_OFN17_gl_rom_n_16, A2 => gl_rom_rom_526(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_527(0), ZN => gl_rom_n_314);
  gl_rom_g36366 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_524(0), B1 => FE_OFN11_gl_rom_n_19, B2 => gl_rom_rom_522(0), ZN => gl_rom_n_313);
  gl_rom_g36367 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_9(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_13(0), ZN => gl_rom_n_312);
  gl_rom_g36368 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_2(1), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_7(1), ZN => gl_rom_n_311);
  gl_rom_g36369 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_4(1), B1 => FE_OFN17_gl_rom_n_16, B2 => gl_rom_rom_6(1), ZN => gl_rom_n_310);
  gl_rom_g36370 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_780(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_782(0), ZN => gl_rom_n_309);
  gl_rom_g36371 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_8(0), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_11(0), ZN => gl_rom_n_308);
  gl_rom_g36372 : AOI22D0BWP7T port map(A1 => FE_OFN14_gl_rom_n_22, A2 => gl_rom_rom_5(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_3(1), ZN => gl_rom_n_307);
  gl_rom_g36373 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_0(1), B1 => FE_OFN25_gl_rom_n_21, B2 => gl_rom_rom_1(1), ZN => gl_rom_n_306);
  gl_rom_g36374 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_6(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_7(0), ZN => gl_rom_n_305);
  gl_rom_g36375 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_521(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_525(0), ZN => gl_rom_n_304);
  gl_rom_g36376 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_4(0), B1 => FE_OFN11_gl_rom_n_19, B2 => gl_rom_rom_2(0), ZN => gl_rom_n_303);
  gl_rom_g36377 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_908(0), B1 => FE_OFN11_gl_rom_n_19, B2 => gl_rom_rom_906(0), ZN => gl_rom_n_302);
  gl_rom_g36378 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_520(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_523(0), ZN => gl_rom_n_301);
  gl_rom_g36379 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_1(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_5(0), ZN => gl_rom_n_300);
  gl_rom_g36380 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_0(0), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_3(0), ZN => gl_rom_n_299);
  gl_rom_g36381 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_778(0), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_779(0), ZN => gl_rom_n_298);
  gl_rom_g36382 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_513(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_517(0), ZN => gl_rom_n_297);
  gl_rom_g36383 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_516(0), B1 => FE_OFN17_gl_rom_n_16, B2 => gl_rom_rom_518(0), ZN => gl_rom_n_296);
  gl_rom_g36384 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_754(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_759(1), ZN => gl_rom_n_295);
  gl_rom_g36385 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_225(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_231(1), ZN => gl_rom_n_294);
  gl_rom_g36386 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_776(0), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_783(0), ZN => gl_rom_n_293);
  gl_rom_g36387 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_757(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_755(1), ZN => gl_rom_n_292);
  gl_rom_g36388 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_514(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_515(0), ZN => gl_rom_n_291);
  gl_rom_g36389 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_752(1), B1 => FE_OFN25_gl_rom_n_21, B2 => gl_rom_rom_753(1), ZN => gl_rom_n_290);
  gl_rom_g36390 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_970(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_973(0), ZN => gl_rom_n_289);
  gl_rom_g36391 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_905(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_909(0), ZN => gl_rom_n_288);
  gl_rom_g36392 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_726(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_727(1), ZN => gl_rom_n_287);
  gl_rom_g36393 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_512(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_519(0), ZN => gl_rom_n_286);
  gl_rom_g36394 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_724(1), B1 => FE_OFN11_gl_rom_n_19, B2 => gl_rom_rom_722(1), ZN => gl_rom_n_285);
  gl_rom_g36395 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_721(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_725(1), ZN => gl_rom_n_284);
  gl_rom_g36396 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_720(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_723(1), ZN => gl_rom_n_283);
  gl_rom_g36397 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_774(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_775(0), ZN => gl_rom_n_282);
  gl_rom_g36398 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_772(0), B1 => FE_OFN11_gl_rom_n_19, B2 => gl_rom_rom_770(0), ZN => gl_rom_n_281);
  gl_rom_g36399 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_730(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_735(1), ZN => gl_rom_n_280);
  gl_rom_g36400 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_904(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_907(0), ZN => gl_rom_n_279);
  gl_rom_g36401 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_732(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_734(1), ZN => gl_rom_n_278);
  gl_rom_g36402 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_250(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_255(0), ZN => gl_rom_n_277);
  gl_rom_g36403 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_733(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_731(1), ZN => gl_rom_n_276);
  gl_rom_g36404 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_252(0), B1 => FE_OFN21_gl_rom_n_16, B2 => gl_rom_rom_254(0), ZN => gl_rom_n_275);
  gl_rom_g36405 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_728(1), B1 => FE_OFN25_gl_rom_n_21, B2 => gl_rom_rom_729(1), ZN => gl_rom_n_274);
  gl_rom_g36406 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_16, A2 => gl_rom_rom_742(1), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_743(1), ZN => gl_rom_n_273);
  gl_rom_g36407 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_740(1), B1 => FE_OFN11_gl_rom_n_19, B2 => gl_rom_rom_738(1), ZN => gl_rom_n_272);
  gl_rom_g36408 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_1010(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_1011(0), ZN => gl_rom_n_271);
  gl_rom_g36409 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_769(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_773(0), ZN => gl_rom_n_270);
  gl_rom_g36410 : AOI22D0BWP7T port map(A1 => FE_OFN16_gl_rom_n_22, A2 => gl_rom_rom_253(0), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_251(0), ZN => gl_rom_n_269);
  gl_rom_g36411 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_737(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_741(1), ZN => gl_rom_n_268);
  gl_rom_g36412 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_736(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_739(1), ZN => gl_rom_n_267);
  gl_rom_g36413 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_248(0), B1 => FE_OFN27_gl_rom_n_21, B2 => gl_rom_rom_249(0), ZN => gl_rom_n_266);
  gl_rom_g36414 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_972(0), B1 => FE_OFN17_gl_rom_n_16, B2 => gl_rom_rom_974(0), ZN => gl_rom_n_265);
  gl_rom_g36415 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_762(1), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_767(1), ZN => gl_rom_n_264);
  gl_rom_g36416 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_764(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_766(1), ZN => gl_rom_n_263);
  gl_rom_g36417 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_768(0), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_771(0), ZN => gl_rom_n_262);
  gl_rom_g36418 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_233(0), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_237(0), ZN => gl_rom_n_261);
  gl_rom_g36419 : AOI22D0BWP7T port map(A1 => FE_OFN15_gl_rom_n_22, A2 => gl_rom_rom_765(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_763(1), ZN => gl_rom_n_260);
  gl_rom_g36420 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_236(0), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_238(0), ZN => gl_rom_n_259);
  gl_rom_g36421 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_760(1), B1 => FE_OFN25_gl_rom_n_21, B2 => gl_rom_rom_761(1), ZN => gl_rom_n_258);
  gl_rom_g36422 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_968(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_971(0), ZN => gl_rom_n_257);
  gl_rom_g36423 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_745(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_749(1), ZN => gl_rom_n_256);
  gl_rom_g36424 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_748(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_750(1), ZN => gl_rom_n_255);
  gl_rom_g36425 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_234(0), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_235(0), ZN => gl_rom_n_254);
  gl_rom_g36426 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_902(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_903(0), ZN => gl_rom_n_253);
  gl_rom_g36427 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_746(1), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_751(1), ZN => gl_rom_n_252);
  gl_rom_g36428 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_232(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_239(0), ZN => gl_rom_n_251);
  gl_rom_g36429 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_744(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_747(1), ZN => gl_rom_n_250);
  gl_rom_g36430 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_900(0), B1 => FE_OFN11_gl_rom_n_19, B2 => gl_rom_rom_898(0), ZN => gl_rom_n_249);
  gl_rom_g36431 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_713(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_717(1), ZN => gl_rom_n_248);
  gl_rom_g36432 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_716(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_718(1), ZN => gl_rom_n_247);
  gl_rom_g36433 : AOI22D0BWP7T port map(A1 => FE_OFN21_gl_rom_n_16, A2 => gl_rom_rom_246(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_247(0), ZN => gl_rom_n_246);
  gl_rom_g36434 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_714(1), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_719(1), ZN => gl_rom_n_245);
  gl_rom_g36435 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_712(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_715(1), ZN => gl_rom_n_244);
  gl_rom_g36436 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_244(0), B1 => FE_OFN13_gl_rom_n_19, B2 => gl_rom_rom_242(0), ZN => gl_rom_n_243);
  gl_rom_g36437 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_886(0), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_887(0), ZN => gl_rom_n_242);
  gl_rom_g36438 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_710(1), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_711(1), ZN => gl_rom_n_241);
  gl_rom_g36439 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_884(0), B1 => FE_OFN12_gl_rom_n_19, B2 => gl_rom_rom_882(0), ZN => gl_rom_n_240);
  gl_rom_g36440 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_708(1), B1 => FE_OFN11_gl_rom_n_19, B2 => gl_rom_rom_706(1), ZN => gl_rom_n_239);
  gl_rom_g36441 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_241(0), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_245(0), ZN => gl_rom_n_238);
  gl_rom_g36442 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_705(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_709(1), ZN => gl_rom_n_237);
  gl_rom_g36443 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_240(0), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_243(0), ZN => gl_rom_n_236);
  gl_rom_g36444 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_704(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_707(1), ZN => gl_rom_n_235);
  gl_rom_g36445 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_793(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_797(1), ZN => gl_rom_n_234);
  gl_rom_g36446 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_796(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_798(1), ZN => gl_rom_n_233);
  gl_rom_g36447 : AOI22D0BWP7T port map(A1 => FE_OFN21_gl_rom_n_16, A2 => gl_rom_rom_214(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_215(0), ZN => gl_rom_n_232);
  gl_rom_g36448 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_897(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_901(0), ZN => gl_rom_n_231);
  gl_rom_g36449 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_881(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_885(0), ZN => gl_rom_n_230);
  gl_rom_g36450 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_794(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_795(1), ZN => gl_rom_n_229);
  gl_rom_g36451 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_792(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_799(1), ZN => gl_rom_n_228);
  gl_rom_g36452 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_212(0), B1 => FE_OFN13_gl_rom_n_19, B2 => gl_rom_rom_210(0), ZN => gl_rom_n_227);
  gl_rom_g36453 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_880(0), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_883(0), ZN => gl_rom_n_226);
  gl_rom_g36454 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_802(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_807(1), ZN => gl_rom_n_225);
  gl_rom_g36455 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_209(0), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_213(0), ZN => gl_rom_n_224);
  gl_rom_g36456 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_801(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_805(1), ZN => gl_rom_n_223);
  gl_rom_g36457 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_208(0), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_211(0), ZN => gl_rom_n_222);
  gl_rom_g36458 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_804(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_803(1), ZN => gl_rom_n_221);
  gl_rom_g36459 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_800(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_806(1), ZN => gl_rom_n_220);
  gl_rom_g36460 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_896(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_899(0), ZN => gl_rom_n_219);
  gl_rom_g36461 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_817(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_821(1), ZN => gl_rom_n_218);
  gl_rom_g36462 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_820(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_822(1), ZN => gl_rom_n_217);
  gl_rom_g36463 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_217(0), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_221(0), ZN => gl_rom_n_216);
  gl_rom_g36464 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_818(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_819(1), ZN => gl_rom_n_215);
  gl_rom_g36465 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_816(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_823(1), ZN => gl_rom_n_214);
  gl_rom_g36466 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_854(0), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_855(0), ZN => gl_rom_n_213);
  gl_rom_g36467 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_220(0), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_222(0), ZN => gl_rom_n_212);
  gl_rom_g36468 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_852(0), B1 => FE_OFN12_gl_rom_n_19, B2 => gl_rom_rom_850(0), ZN => gl_rom_n_211);
  gl_rom_g36469 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_786(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_791(1), ZN => gl_rom_n_210);
  gl_rom_g36470 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_788(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_790(1), ZN => gl_rom_n_209);
  gl_rom_g36471 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_218(0), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_219(0), ZN => gl_rom_n_208);
  gl_rom_g36472 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_789(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_787(1), ZN => gl_rom_n_207);
  gl_rom_g36473 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_784(1), B1 => FE_OFN26_gl_rom_n_21, B2 => gl_rom_rom_785(1), ZN => gl_rom_n_206);
  gl_rom_g36474 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_216(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_223(0), ZN => gl_rom_n_205);
  gl_rom_g36475 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_825(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_829(1), ZN => gl_rom_n_204);
  gl_rom_g36476 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_1008(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_1015(0), ZN => gl_rom_n_203);
  gl_rom_g36477 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_849(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_853(0), ZN => gl_rom_n_202);
  gl_rom_g36478 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_828(1), B1 => FE_OFN19_gl_rom_n_16, B2 => gl_rom_rom_830(1), ZN => gl_rom_n_201);
  gl_rom_g36479 : AOI22D0BWP7T port map(A1 => FE_OFN21_gl_rom_n_16, A2 => gl_rom_rom_230(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_231(0), ZN => gl_rom_n_200);
  gl_rom_g36480 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_826(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_827(1), ZN => gl_rom_n_199);
  gl_rom_g36481 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_228(0), B1 => FE_OFN13_gl_rom_n_19, B2 => gl_rom_rom_226(0), ZN => gl_rom_n_198);
  gl_rom_g36482 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_824(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_831(1), ZN => gl_rom_n_197);
  gl_rom_g36483 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_1016(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_1017(0), ZN => gl_rom_n_196);
  gl_rom_g36484 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_16, A2 => gl_rom_rom_814(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_815(1), ZN => gl_rom_n_195);
  gl_rom_g36485 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_848(0), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_851(0), ZN => gl_rom_n_194);
  gl_rom_g36486 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_225(0), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_229(0), ZN => gl_rom_n_193);
  gl_rom_g36487 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_812(1), B1 => FE_OFN11_gl_rom_n_19, B2 => gl_rom_rom_810(1), ZN => gl_rom_n_192);
  gl_rom_g36488 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_961(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_967(0), ZN => gl_rom_n_191);
  gl_rom_g36489 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_809(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_813(1), ZN => gl_rom_n_190);
  gl_rom_g36490 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_224(0), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_227(0), ZN => gl_rom_n_189);
  gl_rom_g36491 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_808(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_811(1), ZN => gl_rom_n_188);
  gl_rom_g36492 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_777(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_783(1), ZN => gl_rom_n_187);
  gl_rom_g36493 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_778(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_781(1), ZN => gl_rom_n_186);
  gl_rom_g36494 : AOI22D0BWP7T port map(A1 => FE_OFN21_gl_rom_n_16, A2 => gl_rom_rom_206(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_207(0), ZN => gl_rom_n_185);
  gl_rom_g36495 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_780(1), B1 => FE_OFN19_gl_rom_n_16, B2 => gl_rom_rom_782(1), ZN => gl_rom_n_184);
  gl_rom_g36496 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_857(0), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_863(0), ZN => gl_rom_n_183);
  gl_rom_g36497 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_776(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_779(1), ZN => gl_rom_n_182);
  gl_rom_g36498 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_204(0), B1 => FE_OFN13_gl_rom_n_19, B2 => gl_rom_rom_202(0), ZN => gl_rom_n_181);
  gl_rom_g36499 : AOI22D0BWP7T port map(A1 => FE_OFN17_gl_rom_n_16, A2 => gl_rom_rom_766(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_767(0), ZN => gl_rom_n_180);
  gl_rom_g36500 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_769(1), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_775(1), ZN => gl_rom_n_179);
  gl_rom_g36501 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_770(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_773(1), ZN => gl_rom_n_178);
  gl_rom_g36502 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_201(0), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_205(0), ZN => gl_rom_n_177);
  gl_rom_g36503 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_772(1), B1 => FE_OFN19_gl_rom_n_16, B2 => gl_rom_rom_774(1), ZN => gl_rom_n_176);
  gl_rom_g36504 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_200(0), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_203(0), ZN => gl_rom_n_175);
  gl_rom_g36505 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_20, A2 => gl_rom_rom_768(1), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_771(1), ZN => gl_rom_n_174);
  gl_rom_g36506 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_858(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_861(0), ZN => gl_rom_n_173);
  gl_rom_g36507 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_962(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_965(0), ZN => gl_rom_n_172);
  gl_rom_g36508 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_764(0), B1 => gl_rom_n_19, B2 => gl_rom_rom_762(0), ZN => gl_rom_n_171);
  gl_rom_g36509 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_890(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_895(1), ZN => gl_rom_n_170);
  gl_rom_g36510 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_193(0), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_197(0), ZN => gl_rom_n_169);
  gl_rom_g36511 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_892(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_894(1), ZN => gl_rom_n_168);
  gl_rom_g36512 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_860(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_862(0), ZN => gl_rom_n_167);
  gl_rom_g36513 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_196(0), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_198(0), ZN => gl_rom_n_166);
  gl_rom_g36514 : AOI22D0BWP7T port map(A1 => FE_OFN16_gl_rom_n_22, A2 => gl_rom_rom_893(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_891(1), ZN => gl_rom_n_165);
  gl_rom_g36515 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_888(1), B1 => FE_OFN27_gl_rom_n_21, B2 => gl_rom_rom_889(1), ZN => gl_rom_n_164);
  gl_rom_g36516 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_856(0), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_859(0), ZN => gl_rom_n_163);
  gl_rom_g36517 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_194(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_199(0), ZN => gl_rom_n_162);
  gl_rom_g36518 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_874(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_879(1), ZN => gl_rom_n_161);
  gl_rom_g36519 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_876(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_878(1), ZN => gl_rom_n_160);
  gl_rom_g36520 : AOI22D0BWP7T port map(A1 => FE_OFN16_gl_rom_n_22, A2 => gl_rom_rom_877(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_875(1), ZN => gl_rom_n_159);
  gl_rom_g36521 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_872(1), B1 => FE_OFN27_gl_rom_n_21, B2 => gl_rom_rom_873(1), ZN => gl_rom_n_158);
  gl_rom_g36522 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_192(0), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_195(0), ZN => gl_rom_n_157);
  gl_rom_g36523 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_857(1), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_861(1), ZN => gl_rom_n_156);
  gl_rom_g36524 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_761(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_765(0), ZN => gl_rom_n_155);
  gl_rom_g36525 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_860(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_862(1), ZN => gl_rom_n_154);
  gl_rom_g36526 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_870(0), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_871(0), ZN => gl_rom_n_153);
  gl_rom_g36527 : AOI22D0BWP7T port map(A1 => FE_OFN21_gl_rom_n_16, A2 => gl_rom_rom_286(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_287(0), ZN => gl_rom_n_152);
  gl_rom_g36528 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_858(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_863(1), ZN => gl_rom_n_151);
  gl_rom_g36529 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_284(0), B1 => FE_OFN13_gl_rom_n_19, B2 => gl_rom_rom_282(0), ZN => gl_rom_n_150);
  gl_rom_g36530 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_856(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_859(1), ZN => gl_rom_n_149);
  gl_rom_g36531 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_866(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_871(1), ZN => gl_rom_n_148);
  gl_rom_g36532 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_868(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_870(1), ZN => gl_rom_n_147);
  gl_rom_g36533 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_868(0), B1 => FE_OFN12_gl_rom_n_19, B2 => gl_rom_rom_866(0), ZN => gl_rom_n_146);
  gl_rom_g36534 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_281(0), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_285(0), ZN => gl_rom_n_145);
  gl_rom_g36535 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_964(0), B1 => FE_OFN17_gl_rom_n_16, B2 => gl_rom_rom_966(0), ZN => gl_rom_n_144);
  gl_rom_g36536 : AOI22D0BWP7T port map(A1 => FE_OFN16_gl_rom_n_22, A2 => gl_rom_rom_869(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_867(1), ZN => gl_rom_n_143);
  gl_rom_g36537 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_864(1), B1 => FE_OFN27_gl_rom_n_21, B2 => gl_rom_rom_865(1), ZN => gl_rom_n_142);
  gl_rom_g36538 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_280(0), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_283(0), ZN => gl_rom_n_141);
  gl_rom_g36539 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_760(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_763(0), ZN => gl_rom_n_140);
  gl_rom_g36540 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_882(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_887(1), ZN => gl_rom_n_139);
  gl_rom_g36541 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_884(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_886(1), ZN => gl_rom_n_138);
  gl_rom_g36542 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_21, A2 => gl_rom_rom_865(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_869(0), ZN => gl_rom_n_137);
  gl_rom_g36543 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_289(0), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_293(0), ZN => gl_rom_n_136);
  gl_rom_g36544 : AOI22D0BWP7T port map(A1 => FE_OFN16_gl_rom_n_22, A2 => gl_rom_rom_885(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_883(1), ZN => gl_rom_n_135);
  gl_rom_g36545 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_292(0), B1 => FE_OFN21_gl_rom_n_16, B2 => gl_rom_rom_294(0), ZN => gl_rom_n_134);
  gl_rom_g36546 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_880(1), B1 => FE_OFN27_gl_rom_n_21, B2 => gl_rom_rom_881(1), ZN => gl_rom_n_133);
  gl_rom_g36547 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_864(0), B1 => FE_OFN6_gl_rom_n_15, B2 => gl_rom_rom_867(0), ZN => gl_rom_n_132);
  gl_rom_g36548 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_850(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_855(1), ZN => gl_rom_n_131);
  gl_rom_g36549 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_290(0), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_291(0), ZN => gl_rom_n_130);
  gl_rom_g36550 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_852(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_854(1), ZN => gl_rom_n_129);
  gl_rom_g36551 : AOI22D0BWP7T port map(A1 => FE_OFN16_gl_rom_n_22, A2 => gl_rom_rom_853(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_851(1), ZN => gl_rom_n_128);
  gl_rom_g36552 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_288(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_295(0), ZN => gl_rom_n_127);
  gl_rom_g36553 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_848(1), B1 => FE_OFN27_gl_rom_n_21, B2 => gl_rom_rom_849(1), ZN => gl_rom_n_126);
  gl_rom_g36554 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_841(1), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_845(1), ZN => gl_rom_n_125);
  gl_rom_g36555 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_844(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_846(1), ZN => gl_rom_n_124);
  gl_rom_g36556 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_305(0), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_309(0), ZN => gl_rom_n_123);
  gl_rom_g36557 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_889(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_893(0), ZN => gl_rom_n_122);
  gl_rom_g36558 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_842(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_843(1), ZN => gl_rom_n_121);
  gl_rom_g36559 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_840(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_847(1), ZN => gl_rom_n_120);
  gl_rom_g36560 : AOI22D0BWP7T port map(A1 => FE_OFN17_gl_rom_n_16, A2 => gl_rom_rom_750(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_751(0), ZN => gl_rom_n_119);
  gl_rom_g36561 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_308(0), B1 => FE_OFN21_gl_rom_n_16, B2 => gl_rom_rom_310(0), ZN => gl_rom_n_118);
  gl_rom_g36562 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_834(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_839(1), ZN => gl_rom_n_117);
  gl_rom_g36563 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_960(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_963(0), ZN => gl_rom_n_116);
  gl_rom_g36564 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_836(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_838(1), ZN => gl_rom_n_115);
  gl_rom_g36565 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_892(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_894(0), ZN => gl_rom_n_114);
  gl_rom_g36566 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_306(0), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_307(0), ZN => gl_rom_n_113);
  gl_rom_g36567 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_304(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_311(0), ZN => gl_rom_n_112);
  gl_rom_g36568 : AOI22D0BWP7T port map(A1 => FE_OFN16_gl_rom_n_22, A2 => gl_rom_rom_837(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_835(1), ZN => gl_rom_n_111);
  gl_rom_g36569 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_832(1), B1 => FE_OFN27_gl_rom_n_21, B2 => gl_rom_rom_833(1), ZN => gl_rom_n_110);
  gl_rom_g36570 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_748(0), B1 => gl_rom_n_19, B2 => gl_rom_rom_746(0), ZN => gl_rom_n_109);
  gl_rom_g36571 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_634(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_639(1), ZN => gl_rom_n_108);
  gl_rom_g36572 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_274(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_279(0), ZN => gl_rom_n_107);
  gl_rom_g36573 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_636(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_638(1), ZN => gl_rom_n_106);
  gl_rom_g36574 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_890(0), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_891(0), ZN => gl_rom_n_105);
  gl_rom_g36575 : AOI22D0BWP7T port map(A1 => FE_OFN16_gl_rom_n_22, A2 => gl_rom_rom_637(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_635(1), ZN => gl_rom_n_104);
  gl_rom_g36576 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_632(1), B1 => FE_OFN27_gl_rom_n_21, B2 => gl_rom_rom_633(1), ZN => gl_rom_n_103);
  gl_rom_g36577 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_276(0), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_278(0), ZN => gl_rom_n_102);
  gl_rom_g36578 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_888(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_895(0), ZN => gl_rom_n_101);
  gl_rom_g36579 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_618(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_623(1), ZN => gl_rom_n_100);
  gl_rom_g36580 : AOI22D0BWP7T port map(A1 => FE_OFN16_gl_rom_n_22, A2 => gl_rom_rom_277(0), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_275(0), ZN => gl_rom_n_99);
  gl_rom_g36581 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_620(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_622(1), ZN => gl_rom_n_98);
  gl_rom_g36582 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_272(0), B1 => FE_OFN27_gl_rom_n_21, B2 => gl_rom_rom_273(0), ZN => gl_rom_n_97);
  gl_rom_g36583 : AOI22D0BWP7T port map(A1 => FE_OFN16_gl_rom_n_22, A2 => gl_rom_rom_621(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_619(1), ZN => gl_rom_n_96);
  gl_rom_g36584 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_616(1), B1 => FE_OFN27_gl_rom_n_21, B2 => gl_rom_rom_617(1), ZN => gl_rom_n_95);
  gl_rom_g36585 : AOI22D0BWP7T port map(A1 => FE_OFN17_gl_rom_n_16, A2 => gl_rom_rom_982(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_983(0), ZN => gl_rom_n_94);
  gl_rom_g36586 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_601(1), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_605(1), ZN => gl_rom_n_93);
  gl_rom_g36587 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_745(0), B1 => FE_OFN14_gl_rom_n_22, B2 => gl_rom_rom_749(0), ZN => gl_rom_n_92);
  gl_rom_g36588 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_604(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_606(1), ZN => gl_rom_n_91);
  gl_rom_g36589 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_16, A2 => gl_rom_rom_318(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_319(0), ZN => gl_rom_n_90);
  gl_rom_g36590 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_873(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_877(0), ZN => gl_rom_n_89);
  gl_rom_g36591 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_602(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_603(1), ZN => gl_rom_n_88);
  gl_rom_g36592 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_600(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_607(1), ZN => gl_rom_n_87);
  gl_rom_g36593 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_316(0), B1 => FE_OFN13_gl_rom_n_19, B2 => gl_rom_rom_314(0), ZN => gl_rom_n_86);
  gl_rom_g36594 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_876(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_878(0), ZN => gl_rom_n_85);
  gl_rom_g36595 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_609(1), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_613(1), ZN => gl_rom_n_84);
  gl_rom_g36596 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_612(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_614(1), ZN => gl_rom_n_83);
  gl_rom_g36597 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_313(0), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_317(0), ZN => gl_rom_n_82);
  gl_rom_g36598 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_610(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_611(1), ZN => gl_rom_n_81);
  gl_rom_g36599 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_608(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_615(1), ZN => gl_rom_n_80);
  gl_rom_g36600 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_312(0), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_315(0), ZN => gl_rom_n_79);
  gl_rom_g36601 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_1018(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_1023(0), ZN => gl_rom_n_78);
  gl_rom_g36602 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_626(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_631(1), ZN => gl_rom_n_77);
  gl_rom_g36603 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_744(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_747(0), ZN => gl_rom_n_76);
  gl_rom_g36604 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_19, A2 => gl_rom_rom_874(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_879(0), ZN => gl_rom_n_75);
  gl_rom_g36605 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_625(1), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_629(1), ZN => gl_rom_n_74);
  gl_rom_g36606 : AOI22D0BWP7T port map(A1 => FE_OFN21_gl_rom_n_16, A2 => gl_rom_rom_302(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_303(0), ZN => gl_rom_n_73);
  gl_rom_g36607 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_980(0), B1 => gl_rom_n_19, B2 => gl_rom_rom_978(0), ZN => gl_rom_n_72);
  gl_rom_g36608 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_628(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_627(1), ZN => gl_rom_n_71);
  gl_rom_g36609 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_300(0), B1 => FE_OFN13_gl_rom_n_19, B2 => gl_rom_rom_298(0), ZN => gl_rom_n_70);
  gl_rom_g36610 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_624(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_630(1), ZN => gl_rom_n_69);
  gl_rom_g36611 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_20, A2 => gl_rom_rom_872(0), B1 => FE_OFN5_gl_rom_n_15, B2 => gl_rom_rom_875(0), ZN => gl_rom_n_68);
  gl_rom_g36612 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_594(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_599(1), ZN => gl_rom_n_67);
  gl_rom_g36613 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_596(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_598(1), ZN => gl_rom_n_66);
  gl_rom_g36614 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_297(0), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_301(0), ZN => gl_rom_n_65);
  gl_rom_g36615 : AOI22D0BWP7T port map(A1 => FE_OFN16_gl_rom_n_22, A2 => gl_rom_rom_597(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_595(1), ZN => gl_rom_n_64);
  gl_rom_g36616 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_296(0), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_299(0), ZN => gl_rom_n_63);
  gl_rom_g36617 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_592(1), B1 => FE_OFN27_gl_rom_n_21, B2 => gl_rom_rom_593(1), ZN => gl_rom_n_62);
  gl_rom_g36618 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_585(1), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_589(1), ZN => gl_rom_n_61);
  gl_rom_g36619 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_588(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_590(1), ZN => gl_rom_n_60);
  gl_rom_g36620 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_265(0), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_269(0), ZN => gl_rom_n_59);
  gl_rom_g36621 : AOI22D0BWP7T port map(A1 => FE_OFN17_gl_rom_n_16, A2 => gl_rom_rom_758(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_759(0), ZN => gl_rom_n_58);
  gl_rom_g36622 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_846(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_847(0), ZN => gl_rom_n_57);
  gl_rom_g36623 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_586(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_591(1), ZN => gl_rom_n_56);
  gl_rom_g36624 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_268(0), B1 => FE_OFN21_gl_rom_n_16, B2 => gl_rom_rom_270(0), ZN => gl_rom_n_55);
  gl_rom_g36625 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_584(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_587(1), ZN => gl_rom_n_54);
  gl_rom_g36626 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_21, A2 => gl_rom_rom_577(1), B1 => FE_OFN16_gl_rom_n_22, B2 => gl_rom_rom_581(1), ZN => gl_rom_n_53);
  gl_rom_g36627 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_266(0), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_267(0), ZN => gl_rom_n_52);
  gl_rom_g36628 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_580(1), B1 => FE_OFN20_gl_rom_n_16, B2 => gl_rom_rom_582(1), ZN => gl_rom_n_51);
  gl_rom_g36629 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_18, A2 => gl_rom_rom_844(0), B1 => FE_OFN12_gl_rom_n_19, B2 => gl_rom_rom_842(0), ZN => gl_rom_n_50);
  gl_rom_g36630 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_19, A2 => gl_rom_rom_578(1), B1 => FE_OFN7_gl_rom_n_15, B2 => gl_rom_rom_579(1), ZN => gl_rom_n_49);
  gl_rom_g36631 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_576(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_583(1), ZN => gl_rom_n_48);
  gl_rom_g36632 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_20, A2 => gl_rom_rom_264(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_271(0), ZN => gl_rom_n_47);
  gl_rom_g36633 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_950(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_951(0), ZN => gl_rom_n_46);
  gl_rom_g36634 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_756(0), B1 => gl_rom_n_19, B2 => gl_rom_rom_754(0), ZN => gl_rom_n_45);
  gl_rom_g36635 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_21, A2 => gl_rom_rom_1017(1), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_1023(1), ZN => gl_rom_n_44);
  gl_rom_g36636 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_841(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_845(0), ZN => gl_rom_n_43);
  gl_rom_g36637 : AOI22D0BWP7T port map(A1 => FE_OFN21_gl_rom_n_16, A2 => gl_rom_rom_262(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_263(0), ZN => gl_rom_n_42);
  gl_rom_g36638 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_19, A2 => gl_rom_rom_1018(1), B1 => FE_OFN15_gl_rom_n_22, B2 => gl_rom_rom_1021(1), ZN => gl_rom_n_41);
  gl_rom_g36639 : AOI22D0BWP7T port map(A1 => FE_OFN30_gl_rom_n_18, A2 => gl_rom_rom_260(0), B1 => FE_OFN13_gl_rom_n_19, B2 => gl_rom_rom_258(0), ZN => gl_rom_n_40);
  gl_rom_g36640 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_18, A2 => gl_rom_rom_1020(1), B1 => FE_OFN19_gl_rom_n_16, B2 => gl_rom_rom_1022(1), ZN => gl_rom_n_39);
  gl_rom_g36641 : NR2D1BWP7T port map(A1 => gl_rom_n_4, A2 => gl_sig_e(8), ZN => gl_rom_n_38);
  gl_rom_g36642 : INR2D1BWP7T port map(A1 => gl_sig_e(8), B1 => gl_rom_n_1, ZN => gl_rom_n_37);
  gl_rom_g36643 : NR2D1BWP7T port map(A1 => gl_rom_n_9, A2 => gl_sig_e(8), ZN => gl_rom_n_36);
  gl_rom_g36644 : NR2D1BWP7T port map(A1 => gl_rom_n_1, A2 => gl_sig_e(8), ZN => gl_rom_n_35);
  gl_rom_g36645 : INR2D1BWP7T port map(A1 => gl_sig_e(8), B1 => gl_rom_n_4, ZN => gl_rom_n_34);
  gl_rom_g36646 : AN2D1BWP7T port map(A1 => gl_rom_n_10, A2 => gl_sig_e(8), Z => gl_rom_n_33);
  gl_rom_g36647 : INR2D1BWP7T port map(A1 => gl_rom_n_10, B1 => gl_sig_e(8), ZN => gl_rom_n_32);
  gl_rom_g36648 : INR2D1BWP7T port map(A1 => gl_sig_e(8), B1 => gl_rom_n_9, ZN => gl_rom_n_31);
  gl_rom_g36649 : AN2D1BWP7T port map(A1 => gl_rom_n_6, A2 => gl_sig_e(5), Z => gl_rom_n_30);
  gl_rom_g36650 : NR2XD1BWP7T port map(A1 => gl_rom_n_13, A2 => gl_sig_e(5), ZN => gl_rom_n_29);
  gl_rom_g36651 : INR2D2BWP7T port map(A1 => gl_sig_e(5), B1 => gl_rom_n_3, ZN => gl_rom_n_28);
  gl_rom_g36652 : NR2XD1BWP7T port map(A1 => gl_rom_n_3, A2 => gl_sig_e(5), ZN => gl_rom_n_27);
  gl_rom_g36653 : AN2D1BWP7T port map(A1 => gl_rom_n_8, A2 => gl_sig_e(5), Z => gl_rom_n_26);
  gl_rom_g36654 : AN2D1BWP7T port map(A1 => gl_rom_n_14, A2 => gl_sig_e(5), Z => gl_rom_n_25);
  gl_rom_g36655 : INR2D2BWP7T port map(A1 => gl_rom_n_8, B1 => gl_sig_e(5), ZN => gl_rom_n_24);
  gl_rom_g36656 : NR2XD1BWP7T port map(A1 => gl_rom_n_7, A2 => gl_sig_e(5), ZN => gl_rom_n_23);
  gl_rom_g36657 : AN2D2BWP7T port map(A1 => gl_rom_n_2, A2 => gl_sig_e(2), Z => gl_rom_n_22);
  gl_rom_g36658 : AN2D1BWP7T port map(A1 => gl_rom_n_2, A2 => gl_rom_n_0, Z => gl_rom_n_21);
  gl_rom_g36659 : AN2D2BWP7T port map(A1 => gl_rom_n_5, A2 => gl_rom_n_0, Z => gl_rom_n_20);
  gl_rom_g36660 : AN2D1BWP7T port map(A1 => gl_rom_n_11, A2 => gl_rom_n_0, Z => gl_rom_n_19);
  gl_rom_g36661 : AN2D2BWP7T port map(A1 => gl_rom_n_5, A2 => gl_sig_e(2), Z => gl_rom_n_18);
  gl_rom_g36662 : AN2D2BWP7T port map(A1 => gl_rom_n_12, A2 => gl_sig_e(2), Z => gl_rom_n_17);
  gl_rom_g36663 : AN2D2BWP7T port map(A1 => gl_rom_n_11, A2 => gl_sig_e(2), Z => gl_rom_n_16);
  gl_rom_g36664 : AN2D1BWP7T port map(A1 => gl_rom_n_12, A2 => gl_rom_n_0, Z => gl_rom_n_15);
  gl_rom_g36665 : INVD0BWP7T port map(I => gl_rom_n_13, ZN => gl_rom_n_14);
  gl_rom_g36666 : IND2D1BWP7T port map(A1 => gl_sig_e(4), B1 => gl_sig_e(3), ZN => gl_rom_n_13);
  gl_rom_g36667 : AN2D1BWP7T port map(A1 => gl_sig_e(1), A2 => gl_sig_e(0), Z => gl_rom_n_12);
  gl_rom_g36668 : INR2D1BWP7T port map(A1 => gl_sig_e(1), B1 => gl_sig_e(0), ZN => gl_rom_n_11);
  gl_rom_g36669 : NR2D0BWP7T port map(A1 => gl_sig_e(7), A2 => gl_sig_e(6), ZN => gl_rom_n_10);
  gl_rom_g36670 : ND2D1BWP7T port map(A1 => gl_sig_e(7), A2 => gl_sig_e(6), ZN => gl_rom_n_9);
  gl_rom_g36671 : NR2XD0BWP7T port map(A1 => gl_sig_e(4), A2 => gl_sig_e(3), ZN => gl_rom_n_8);
  gl_rom_g36672 : INVD0BWP7T port map(I => gl_rom_n_6, ZN => gl_rom_n_7);
  gl_rom_g36673 : INR2D1BWP7T port map(A1 => gl_sig_e(4), B1 => gl_sig_e(3), ZN => gl_rom_n_6);
  gl_rom_g36674 : NR2D1BWP7T port map(A1 => gl_sig_e(1), A2 => gl_sig_e(0), ZN => gl_rom_n_5);
  gl_rom_g36675 : IND2D1BWP7T port map(A1 => gl_sig_e(7), B1 => gl_sig_e(6), ZN => gl_rom_n_4);
  gl_rom_g36676 : ND2D1BWP7T port map(A1 => gl_sig_e(4), A2 => gl_sig_e(3), ZN => gl_rom_n_3);
  gl_rom_g36677 : INR2D1BWP7T port map(A1 => gl_sig_e(0), B1 => gl_sig_e(1), ZN => gl_rom_n_2);
  gl_rom_g36678 : IND2D1BWP7T port map(A1 => gl_sig_e(6), B1 => gl_sig_e(7), ZN => gl_rom_n_1);
  gl_rom_g36679 : INVD1BWP7T port map(I => gl_sig_e(2), ZN => gl_rom_n_0);
  gl_ram_g8810 : OAI211D1BWP7T port map(A1 => gl_ram_n_1078, A2 => gl_ram_n_1106, B => gl_ram_n_1109, C => gl_ram_n_1099, ZN => gl_sig_ram(2));
  gl_ram_g8811 : OAI211D1BWP7T port map(A1 => gl_ram_n_1078, A2 => gl_ram_n_1104, B => gl_ram_n_1108, C => gl_ram_n_1102, ZN => gl_sig_ram(0));
  gl_ram_g8812 : OAI211D1BWP7T port map(A1 => gl_ram_n_1078, A2 => gl_ram_n_1105, B => gl_ram_n_1107, C => gl_ram_n_1098, ZN => gl_sig_ram(1));
  gl_ram_g8813 : AOI22D0BWP7T port map(A1 => gl_ram_n_1100, A2 => gl_ram_n_1078, B1 => gl_ram_n_1045, B2 => gl_ram_n_1096, ZN => gl_ram_n_1109);
  gl_ram_g8814 : AOI22D0BWP7T port map(A1 => gl_ram_n_1103, A2 => gl_ram_n_1078, B1 => gl_ram_n_1036, B2 => gl_ram_n_1096, ZN => gl_ram_n_1108);
  gl_ram_g8815 : AOI22D0BWP7T port map(A1 => gl_ram_n_1101, A2 => gl_ram_n_1078, B1 => gl_ram_n_1027, B2 => gl_ram_n_1096, ZN => gl_ram_n_1107);
  gl_ram_g8816 : AOI221D0BWP7T port map(A1 => FE_OCPN239_gl_ram_ram_86_2, A2 => gl_ram_n_1079, B1 => FE_OCPN219_gl_ram_ram_87_2, B2 => gl_ram_n_818, C => gl_ram_n_1092, ZN => gl_ram_n_1106);
  gl_ram_g8817 : AOI221D0BWP7T port map(A1 => FE_OCPN146_gl_ram_ram_86_1, A2 => gl_ram_n_1079, B1 => FE_OCPN144_gl_ram_ram_87_1, B2 => gl_ram_n_818, C => gl_ram_n_1090, ZN => gl_ram_n_1105);
  gl_ram_g8818 : AOI221D0BWP7T port map(A1 => gl_ram_ram_86(0), A2 => gl_ram_n_1079, B1 => gl_ram_ram_87(0), B2 => gl_ram_n_818, C => gl_ram_n_1091, ZN => gl_ram_n_1104);
  gl_ram_g8819 : ND4D0BWP7T port map(A1 => gl_ram_n_1080, A2 => gl_ram_n_1088, A3 => gl_ram_n_1087, A4 => gl_ram_n_1083, ZN => gl_ram_n_1103);
  gl_ram_g8820 : AOI22D0BWP7T port map(A1 => gl_ram_n_1040, A2 => gl_ram_n_1097, B1 => gl_ram_n_1042, B2 => gl_ram_n_1095, ZN => gl_ram_n_1102);
  gl_ram_g8821 : ND4D0BWP7T port map(A1 => gl_ram_n_1089, A2 => gl_ram_n_1093, A3 => gl_ram_n_1081, A4 => gl_ram_n_1085, ZN => gl_ram_n_1101);
  gl_ram_g8822 : ND4D0BWP7T port map(A1 => gl_ram_n_1094, A2 => gl_ram_n_1086, A3 => gl_ram_n_1082, A4 => gl_ram_n_1084, ZN => gl_ram_n_1100);
  gl_ram_g8823 : AOI22D0BWP7T port map(A1 => gl_ram_n_1039, A2 => gl_ram_n_1097, B1 => gl_ram_n_1056, B2 => gl_ram_n_1095, ZN => gl_ram_n_1099);
  gl_ram_g8824 : AOI22D0BWP7T port map(A1 => gl_ram_n_1034, A2 => gl_ram_n_1097, B1 => gl_ram_n_1037, B2 => gl_ram_n_1095, ZN => gl_ram_n_1098);
  gl_ram_g8825 : AOI22D0BWP7T port map(A1 => gl_ram_n_1031, A2 => gl_ram_n_1071, B1 => gl_ram_n_1038, B2 => gl_ram_n_1072, ZN => gl_ram_n_1094);
  gl_ram_g8826 : AOI22D0BWP7T port map(A1 => gl_ram_n_1051, A2 => gl_ram_n_1074, B1 => gl_ram_n_1052, B2 => gl_ram_n_1071, ZN => gl_ram_n_1093);
  gl_ram_g8827 : MOAI22D0BWP7T port map(A1 => gl_ram_n_1023, A2 => gl_ram_n_1075, B1 => gl_ram_n_1050, B2 => gl_ram_n_1073, ZN => gl_ram_n_1092);
  gl_ram_g8828 : MOAI22D0BWP7T port map(A1 => gl_ram_n_1022, A2 => gl_ram_n_1075, B1 => gl_ram_n_1058, B2 => gl_ram_n_1073, ZN => gl_ram_n_1091);
  gl_ram_g8829 : MOAI22D0BWP7T port map(A1 => gl_ram_n_1021, A2 => gl_ram_n_1075, B1 => gl_ram_n_1057, B2 => gl_ram_n_1073, ZN => gl_ram_n_1090);
  gl_ram_g8830 : AOI22D0BWP7T port map(A1 => gl_ram_n_1054, A2 => gl_ram_n_1072, B1 => gl_ram_n_1055, B2 => gl_ram_n_1077, ZN => gl_ram_n_1089);
  gl_ram_g8831 : NR2D1BWP7T port map(A1 => gl_ram_n_1078, A2 => gl_ram_n_1069, ZN => gl_ram_n_1097);
  gl_ram_g8832 : INR2D1BWP7T port map(A1 => gl_ram_n_1070, B1 => gl_ram_n_1078, ZN => gl_ram_n_1096);
  gl_ram_g8833 : INR2D1BWP7T port map(A1 => gl_ram_n_1076, B1 => gl_ram_n_1078, ZN => gl_ram_n_1095);
  gl_ram_g8834 : AOI22D0BWP7T port map(A1 => gl_ram_n_1030, A2 => gl_ram_n_1070, B1 => gl_ram_n_1041, B2 => gl_ram_n_1076, ZN => gl_ram_n_1088);
  gl_ram_g8835 : AOI22D0BWP7T port map(A1 => gl_ram_n_1028, A2 => gl_ram_n_1071, B1 => gl_ram_n_1029, B2 => gl_ram_n_1072, ZN => gl_ram_n_1087);
  gl_ram_g8836 : AOI22D0BWP7T port map(A1 => gl_ram_n_1053, A2 => gl_ram_n_1074, B1 => gl_ram_n_1024, B2 => gl_ram_n_1077, ZN => gl_ram_n_1086);
  gl_ram_g8837 : MAOI22D0BWP7T port map(A1 => gl_ram_n_1046, A2 => gl_ram_n_1073, B1 => gl_ram_n_1044, B2 => gl_ram_n_1069, ZN => gl_ram_n_1085);
  gl_ram_g8838 : MAOI22D0BWP7T port map(A1 => gl_ram_n_1043, A2 => gl_ram_n_1073, B1 => gl_ram_n_1032, B2 => gl_ram_n_1069, ZN => gl_ram_n_1084);
  gl_ram_g8839 : MAOI22D0BWP7T port map(A1 => gl_ram_n_1026, A2 => gl_ram_n_1073, B1 => gl_ram_n_1025, B2 => gl_ram_n_1069, ZN => gl_ram_n_1083);
  gl_ram_g8840 : AOI22D0BWP7T port map(A1 => gl_ram_n_1047, A2 => gl_ram_n_1070, B1 => gl_ram_n_1059, B2 => gl_ram_n_1076, ZN => gl_ram_n_1082);
  gl_ram_g8841 : AOI22D0BWP7T port map(A1 => gl_ram_n_1048, A2 => gl_ram_n_1070, B1 => gl_ram_n_1049, B2 => gl_ram_n_1076, ZN => gl_ram_n_1081);
  gl_ram_g8842 : AOI22D0BWP7T port map(A1 => gl_ram_n_1033, A2 => gl_ram_n_1074, B1 => gl_ram_n_1035, B2 => gl_ram_n_1077, ZN => gl_ram_n_1080);
  gl_ram_g8843 : AN2D1BWP7T port map(A1 => gl_ram_n_1073, A2 => gl_ram_n_873, Z => gl_ram_n_1079);
  gl_ram_g8845 : XNR2D1BWP7T port map(A1 => gl_ram_n_1067, A2 => gl_sig_y(3), ZN => gl_ram_n_1078);
  gl_ram_g8846 : INVD1BWP7T port map(I => gl_ram_n_1075, ZN => gl_ram_n_1074);
  gl_ram_g8847 : INR2D1BWP7T port map(A1 => gl_ram_n_1068, B1 => gl_ram_n_1065, ZN => gl_ram_n_1077);
  gl_ram_g8848 : NR2D1BWP7T port map(A1 => gl_ram_n_1068, A2 => gl_ram_n_1065, ZN => gl_ram_n_1076);
  gl_ram_g8849 : ND2D1BWP7T port map(A1 => gl_ram_n_1068, A2 => gl_ram_n_1062, ZN => gl_ram_n_1075);
  gl_ram_g8850 : NR2D1BWP7T port map(A1 => gl_ram_n_1068, A2 => gl_ram_n_1066, ZN => gl_ram_n_1073);
  gl_ram_g8851 : INR2D1BWP7T port map(A1 => gl_ram_n_1068, B1 => gl_ram_n_1066, ZN => gl_ram_n_1072);
  gl_ram_g8852 : AN2D1BWP7T port map(A1 => gl_ram_n_1068, A2 => gl_ram_n_1063, Z => gl_ram_n_1071);
  gl_ram_g8853 : NR2D1BWP7T port map(A1 => gl_ram_n_1068, A2 => gl_ram_n_1064, ZN => gl_ram_n_1070);
  gl_ram_g8854 : IND2D1BWP7T port map(A1 => gl_ram_n_1068, B1 => gl_ram_n_1062, ZN => gl_ram_n_1069);
  gl_ram_g8855 : FA1D0BWP7T port map(A => gl_ram_n_855, B => gl_sig_y(2), CI => gl_ram_n_1060, CO => gl_ram_n_1067, S => gl_ram_n_1068);
  gl_ram_g8856 : IND2D1BWP7T port map(A1 => gl_ram_n_876, B1 => gl_ram_n_1061, ZN => gl_ram_n_1066);
  gl_ram_g8857 : ND2D1BWP7T port map(A1 => gl_ram_n_1061, A2 => gl_ram_n_876, ZN => gl_ram_n_1065);
  gl_ram_g8858 : INVD0BWP7T port map(I => gl_ram_n_1063, ZN => gl_ram_n_1064);
  gl_ram_g8859 : INR2D1BWP7T port map(A1 => gl_ram_n_876, B1 => gl_ram_n_1061, ZN => gl_ram_n_1063);
  gl_ram_g8860 : NR2D1BWP7T port map(A1 => gl_ram_n_1061, A2 => gl_ram_n_876, ZN => gl_ram_n_1062);
  gl_ram_g8861 : FA1D0BWP7T port map(A => gl_ram_n_856, B => gl_ram_n_857, CI => gl_ram_n_875, CO => gl_ram_n_1060, S => gl_ram_n_1061);
  gl_ram_g8862 : ND4D0BWP7T port map(A1 => gl_ram_n_996, A2 => gl_ram_n_994, A3 => gl_ram_n_988, A4 => gl_ram_n_986, ZN => gl_ram_n_1059);
  gl_ram_g8863 : ND3D0BWP7T port map(A1 => gl_ram_n_946, A2 => gl_ram_n_945, A3 => gl_ram_n_943, ZN => gl_ram_n_1058);
  gl_ram_g8864 : ND3D0BWP7T port map(A1 => gl_ram_n_901, A2 => gl_ram_n_897, A3 => gl_ram_n_893, ZN => gl_ram_n_1057);
  gl_ram_g8865 : ND4D0BWP7T port map(A1 => gl_ram_n_914, A2 => gl_ram_n_910, A3 => gl_ram_n_991, A4 => gl_ram_n_955, ZN => gl_ram_n_1056);
  gl_ram_g8866 : ND4D0BWP7T port map(A1 => gl_ram_n_1019, A2 => gl_ram_n_1018, A3 => gl_ram_n_1016, A4 => gl_ram_n_1015, ZN => gl_ram_n_1055);
  gl_ram_g8867 : ND4D0BWP7T port map(A1 => gl_ram_n_1013, A2 => gl_ram_n_1012, A3 => gl_ram_n_1010, A4 => gl_ram_n_1008, ZN => gl_ram_n_1054);
  gl_ram_g8868 : ND4D0BWP7T port map(A1 => gl_ram_n_1009, A2 => gl_ram_n_1007, A3 => gl_ram_n_1004, A4 => gl_ram_n_1001, ZN => gl_ram_n_1053);
  gl_ram_g8869 : ND4D0BWP7T port map(A1 => gl_ram_n_1006, A2 => gl_ram_n_1005, A3 => gl_ram_n_1003, A4 => gl_ram_n_1002, ZN => gl_ram_n_1052);
  gl_ram_g8870 : ND4D0BWP7T port map(A1 => gl_ram_n_1000, A2 => gl_ram_n_999, A3 => gl_ram_n_998, A4 => gl_ram_n_995, ZN => gl_ram_n_1051);
  gl_ram_g8871 : ND3D0BWP7T port map(A1 => gl_ram_n_997, A2 => gl_ram_n_990, A3 => gl_ram_n_982, ZN => gl_ram_n_1050);
  gl_ram_g8872 : ND4D0BWP7T port map(A1 => gl_ram_n_993, A2 => gl_ram_n_992, A3 => gl_ram_n_989, A4 => gl_ram_n_987, ZN => gl_ram_n_1049);
  gl_ram_g8873 : ND4D0BWP7T port map(A1 => gl_ram_n_985, A2 => gl_ram_n_984, A3 => gl_ram_n_983, A4 => gl_ram_n_981, ZN => gl_ram_n_1048);
  gl_ram_g8874 : ND4D0BWP7T port map(A1 => gl_ram_n_980, A2 => gl_ram_n_979, A3 => gl_ram_n_976, A4 => gl_ram_n_972, ZN => gl_ram_n_1047);
  gl_ram_g8875 : ND4D0BWP7T port map(A1 => gl_ram_n_978, A2 => gl_ram_n_977, A3 => gl_ram_n_975, A4 => gl_ram_n_974, ZN => gl_ram_n_1046);
  gl_ram_g8876 : ND4D0BWP7T port map(A1 => gl_ram_n_973, A2 => gl_ram_n_963, A3 => gl_ram_n_962, A4 => gl_ram_n_954, ZN => gl_ram_n_1045);
  gl_ram_g8877 : AN4D0BWP7T port map(A1 => gl_ram_n_971, A2 => gl_ram_n_970, A3 => gl_ram_n_969, A4 => gl_ram_n_967, Z => gl_ram_n_1044);
  gl_ram_g8878 : ND4D0BWP7T port map(A1 => gl_ram_n_968, A2 => gl_ram_n_966, A3 => gl_ram_n_961, A4 => gl_ram_n_958, ZN => gl_ram_n_1043);
  gl_ram_g8879 : ND4D0BWP7T port map(A1 => gl_ram_n_965, A2 => gl_ram_n_964, A3 => gl_ram_n_960, A4 => gl_ram_n_959, ZN => gl_ram_n_1042);
  gl_ram_g8880 : ND4D0BWP7T port map(A1 => gl_ram_n_917, A2 => gl_ram_n_915, A3 => gl_ram_n_913, A4 => gl_ram_n_911, ZN => gl_ram_n_1041);
  gl_ram_g8881 : ND4D0BWP7T port map(A1 => gl_ram_n_957, A2 => gl_ram_n_956, A3 => gl_ram_n_952, A4 => gl_ram_n_951, ZN => gl_ram_n_1040);
  gl_ram_g8882 : ND4D0BWP7T port map(A1 => gl_ram_n_944, A2 => gl_ram_n_929, A3 => gl_ram_n_918, A4 => gl_ram_n_912, ZN => gl_ram_n_1039);
  gl_ram_g8883 : ND4D0BWP7T port map(A1 => gl_ram_n_939, A2 => gl_ram_n_935, A3 => gl_ram_n_927, A4 => gl_ram_n_921, ZN => gl_ram_n_1038);
  gl_ram_g8884 : ND4D0BWP7T port map(A1 => gl_ram_n_941, A2 => gl_ram_n_938, A3 => gl_ram_n_934, A4 => gl_ram_n_933, ZN => gl_ram_n_1037);
  gl_ram_g8885 : ND4D0BWP7T port map(A1 => gl_ram_n_942, A2 => gl_ram_n_940, A3 => gl_ram_n_937, A4 => gl_ram_n_936, ZN => gl_ram_n_1036);
  gl_ram_g8886 : ND4D0BWP7T port map(A1 => gl_ram_n_932, A2 => gl_ram_n_931, A3 => gl_ram_n_930, A4 => gl_ram_n_928, ZN => gl_ram_n_1035);
  gl_ram_g8887 : ND4D0BWP7T port map(A1 => gl_ram_n_926, A2 => gl_ram_n_923, A3 => gl_ram_n_919, A4 => gl_ram_n_916, ZN => gl_ram_n_1034);
  gl_ram_g8888 : ND4D0BWP7T port map(A1 => gl_ram_n_925, A2 => gl_ram_n_924, A3 => gl_ram_n_922, A4 => gl_ram_n_920, ZN => gl_ram_n_1033);
  gl_ram_g8889 : AN4D0BWP7T port map(A1 => gl_ram_n_953, A2 => gl_ram_n_950, A3 => gl_ram_n_877, A4 => gl_ram_n_947, Z => gl_ram_n_1032);
  gl_ram_g8890 : ND4D0BWP7T port map(A1 => gl_ram_n_908, A2 => gl_ram_n_896, A3 => gl_ram_n_898, A4 => gl_ram_n_891, ZN => gl_ram_n_1031);
  gl_ram_g8891 : ND4D0BWP7T port map(A1 => gl_ram_n_909, A2 => gl_ram_n_907, A3 => gl_ram_n_906, A4 => gl_ram_n_905, ZN => gl_ram_n_1030);
  gl_ram_g8892 : ND4D0BWP7T port map(A1 => gl_ram_n_904, A2 => gl_ram_n_903, A3 => gl_ram_n_900, A4 => gl_ram_n_899, ZN => gl_ram_n_1029);
  gl_ram_g8893 : ND4D0BWP7T port map(A1 => gl_ram_n_895, A2 => gl_ram_n_894, A3 => gl_ram_n_892, A4 => gl_ram_n_890, ZN => gl_ram_n_1028);
  gl_ram_g8894 : ND4D0BWP7T port map(A1 => gl_ram_n_888, A2 => gl_ram_n_886, A3 => gl_ram_n_883, A4 => gl_ram_n_879, ZN => gl_ram_n_1027);
  gl_ram_g8895 : ND4D0BWP7T port map(A1 => gl_ram_n_889, A2 => gl_ram_n_887, A3 => gl_ram_n_885, A4 => gl_ram_n_884, ZN => gl_ram_n_1026);
  gl_ram_g8896 : AN4D0BWP7T port map(A1 => gl_ram_n_882, A2 => gl_ram_n_881, A3 => gl_ram_n_878, A4 => gl_ram_n_948, Z => gl_ram_n_1025);
  gl_ram_g8897 : ND4D0BWP7T port map(A1 => gl_ram_n_880, A2 => gl_ram_n_949, A3 => gl_ram_n_1017, A4 => gl_ram_n_1014, ZN => gl_ram_n_1024);
  gl_ram_g8898 : AOI221D0BWP7T port map(A1 => FE_OCPN38_gl_ram_ram_98_2, A2 => gl_ram_n_868, B1 => gl_ram_ram_97(2), B2 => gl_ram_n_869, C => gl_ram_n_1011, ZN => gl_ram_n_1023);
  gl_ram_g8899 : AOI221D0BWP7T port map(A1 => FE_OCPN36_gl_ram_ram_98_0, A2 => gl_ram_n_868, B1 => gl_ram_ram_97(0), B2 => gl_ram_n_869, C => gl_ram_n_1020, ZN => gl_ram_n_1022);
  gl_ram_g8900 : AOI221D0BWP7T port map(A1 => gl_ram_ram_96(1), A2 => gl_ram_n_867, B1 => FE_OCPN37_gl_ram_ram_97_1, B2 => gl_ram_n_869, C => gl_ram_n_902, ZN => gl_ram_n_1021);
  gl_ram_g8901 : AO22D0BWP7T port map(A1 => gl_ram_ram_99(0), A2 => gl_ram_n_871, B1 => gl_ram_n_867, B2 => gl_ram_ram_96(0), Z => gl_ram_n_1020);
  gl_ram_g8902 : AOI22D0BWP7T port map(A1 => gl_ram_ram_60(1), A2 => gl_ram_n_870, B1 => gl_ram_ram_61(1), B2 => gl_ram_n_872, ZN => gl_ram_n_1019);
  gl_ram_g8903 : AOI22D0BWP7T port map(A1 => gl_ram_ram_62(1), A2 => gl_ram_n_873, B1 => gl_ram_ram_63(1), B2 => gl_ram_n_874, ZN => gl_ram_n_1018);
  gl_ram_g8904 : AOI22D0BWP7T port map(A1 => gl_ram_ram_62(2), A2 => gl_ram_n_873, B1 => gl_ram_ram_63(2), B2 => gl_ram_n_874, ZN => gl_ram_n_1017);
  gl_ram_g8905 : AOI22D0BWP7T port map(A1 => gl_ram_ram_59(1), A2 => gl_ram_n_871, B1 => gl_ram_ram_56(1), B2 => gl_ram_n_867, ZN => gl_ram_n_1016);
  gl_ram_g8906 : AOI22D0BWP7T port map(A1 => gl_ram_ram_58(1), A2 => gl_ram_n_868, B1 => gl_ram_ram_57(1), B2 => gl_ram_n_869, ZN => gl_ram_n_1015);
  gl_ram_g8907 : AOI22D0BWP7T port map(A1 => FE_OCPN159_gl_ram_ram_59_2, A2 => gl_ram_n_871, B1 => gl_ram_ram_56(2), B2 => gl_ram_n_867, ZN => gl_ram_n_1014);
  gl_ram_g8908 : AOI22D0BWP7T port map(A1 => gl_ram_ram_52(1), A2 => gl_ram_n_870, B1 => gl_ram_ram_53(1), B2 => gl_ram_n_872, ZN => gl_ram_n_1013);
  gl_ram_g8909 : AOI22D0BWP7T port map(A1 => FE_OCPN136_gl_ram_ram_51_1, A2 => gl_ram_n_871, B1 => FE_OCPN54_gl_ram_ram_48_1, B2 => gl_ram_n_867, ZN => gl_ram_n_1012);
  gl_ram_g8910 : AO22D0BWP7T port map(A1 => FE_OCPN179_gl_ram_ram_99_2, A2 => gl_ram_n_871, B1 => gl_ram_n_867, B2 => gl_ram_ram_96(2), Z => gl_ram_n_1011);
  gl_ram_g8911 : AOI22D0BWP7T port map(A1 => FE_OCPN184_gl_ram_ram_54_1, A2 => gl_ram_n_873, B1 => FE_OCPN242_gl_ram_ram_55_1, B2 => gl_ram_n_874, ZN => gl_ram_n_1010);
  gl_ram_g8912 : AOI22D0BWP7T port map(A1 => FE_PSN353_gl_ram_ram_36_2, A2 => gl_ram_n_870, B1 => gl_ram_ram_37(2), B2 => gl_ram_n_872, ZN => gl_ram_n_1009);
  gl_ram_g8913 : AOI22D0BWP7T port map(A1 => gl_ram_ram_50(1), A2 => gl_ram_n_868, B1 => gl_ram_ram_49(1), B2 => gl_ram_n_869, ZN => gl_ram_n_1008);
  gl_ram_g8914 : AOI22D0BWP7T port map(A1 => gl_ram_ram_34(2), A2 => gl_ram_n_868, B1 => gl_ram_ram_33(2), B2 => gl_ram_n_869, ZN => gl_ram_n_1007);
  gl_ram_g8915 : AOI22D0BWP7T port map(A1 => gl_ram_ram_44(1), A2 => gl_ram_n_870, B1 => gl_ram_n_872, B2 => gl_ram_ram_45(1), ZN => gl_ram_n_1006);
  gl_ram_g8916 : AOI22D0BWP7T port map(A1 => gl_ram_ram_42(1), A2 => gl_ram_n_868, B1 => FE_OCPN2_gl_ram_ram_41_1, B2 => gl_ram_n_869, ZN => gl_ram_n_1005);
  gl_ram_g8917 : AOI22D0BWP7T port map(A1 => gl_ram_ram_38(2), A2 => gl_ram_n_873, B1 => gl_ram_ram_39(2), B2 => gl_ram_n_874, ZN => gl_ram_n_1004);
  gl_ram_g8918 : AOI22D0BWP7T port map(A1 => gl_ram_ram_46(1), A2 => gl_ram_n_873, B1 => gl_ram_n_874, B2 => FE_OCPN8_gl_ram_ram_47_1, ZN => gl_ram_n_1003);
  gl_ram_g8919 : AOI22D0BWP7T port map(A1 => gl_ram_ram_43(1), A2 => gl_ram_n_871, B1 => FE_OCPN7_gl_ram_ram_40_1, B2 => gl_ram_n_867, ZN => gl_ram_n_1002);
  gl_ram_g8920 : AOI22D0BWP7T port map(A1 => gl_ram_ram_35(2), A2 => gl_ram_n_871, B1 => FE_OCPN77_gl_ram_ram_32_2, B2 => gl_ram_n_867, ZN => gl_ram_n_1001);
  gl_ram_g8921 : AOI22D0BWP7T port map(A1 => gl_ram_ram_36(1), A2 => gl_ram_n_870, B1 => gl_ram_ram_37(1), B2 => gl_ram_n_872, ZN => gl_ram_n_1000);
  gl_ram_g8922 : AOI22D0BWP7T port map(A1 => gl_ram_ram_35(1), A2 => gl_ram_n_871, B1 => FE_OCPN274_gl_ram_ram_32_1, B2 => gl_ram_n_867, ZN => gl_ram_n_999);
  gl_ram_g8923 : AOI22D0BWP7T port map(A1 => gl_ram_ram_38(1), A2 => gl_ram_n_873, B1 => gl_ram_ram_39(1), B2 => gl_ram_n_874, ZN => gl_ram_n_998);
  gl_ram_g8924 : AOI22D0BWP7T port map(A1 => gl_ram_ram_84(2), A2 => gl_ram_n_870, B1 => FE_PSN352_gl_ram_ram_85_2, B2 => gl_ram_n_872, ZN => gl_ram_n_997);
  gl_ram_g8925 : AOI22D0BWP7T port map(A1 => gl_ram_ram_28(2), A2 => gl_ram_n_870, B1 => FE_OCPN244_gl_ram_ram_29_2, B2 => gl_ram_n_872, ZN => gl_ram_n_996);
  gl_ram_g8926 : AOI22D0BWP7T port map(A1 => gl_ram_ram_34(1), A2 => gl_ram_n_868, B1 => FE_OCPN56_gl_ram_ram_33_1, B2 => gl_ram_n_869, ZN => gl_ram_n_995);
  gl_ram_g8927 : AOI22D0BWP7T port map(A1 => gl_ram_ram_30(2), A2 => gl_ram_n_873, B1 => gl_ram_ram_31(2), B2 => gl_ram_n_874, ZN => gl_ram_n_994);
  gl_ram_g8928 : AOI22D0BWP7T port map(A1 => FE_OCPN14_gl_ram_ram_28_1, A2 => gl_ram_n_870, B1 => gl_ram_ram_29(1), B2 => gl_ram_n_872, ZN => gl_ram_n_993);
  gl_ram_g8929 : AOI22D0BWP7T port map(A1 => FE_OCPN6_gl_ram_ram_30_1, A2 => gl_ram_n_873, B1 => gl_ram_ram_31(1), B2 => gl_ram_n_874, ZN => gl_ram_n_992);
  gl_ram_g8930 : AOI22D0BWP7T port map(A1 => gl_ram_ram_94(2), A2 => gl_ram_n_873, B1 => gl_ram_ram_95(2), B2 => gl_ram_n_874, ZN => gl_ram_n_991);
  gl_ram_g8931 : AOI22D0BWP7T port map(A1 => FE_OCPN225_gl_ram_ram_80_2, A2 => gl_ram_n_867, B1 => gl_ram_ram_81(2), B2 => gl_ram_n_869, ZN => gl_ram_n_990);
  gl_ram_g8932 : AOI22D0BWP7T port map(A1 => gl_ram_ram_24(1), A2 => gl_ram_n_867, B1 => FE_OCPN10_gl_ram_ram_25_1, B2 => gl_ram_n_869, ZN => gl_ram_n_989);
  gl_ram_g8933 : AOI22D0BWP7T port map(A1 => gl_ram_ram_27(2), A2 => gl_ram_n_871, B1 => FE_OCPN250_gl_ram_ram_24_2, B2 => gl_ram_n_867, ZN => gl_ram_n_988);
  gl_ram_g8934 : AOI22D0BWP7T port map(A1 => gl_ram_ram_26(1), A2 => gl_ram_n_868, B1 => gl_ram_ram_27(1), B2 => gl_ram_n_871, ZN => gl_ram_n_987);
  gl_ram_g8935 : AOI22D0BWP7T port map(A1 => gl_ram_ram_26(2), A2 => gl_ram_n_868, B1 => FE_OCPN252_gl_ram_ram_25_2, B2 => gl_ram_n_869, ZN => gl_ram_n_986);
  gl_ram_g8936 : AOI22D0BWP7T port map(A1 => FE_OCPN233_gl_ram_ram_12_1, A2 => gl_ram_n_870, B1 => gl_ram_ram_13(1), B2 => gl_ram_n_872, ZN => gl_ram_n_985);
  gl_ram_g8937 : AOI22D0BWP7T port map(A1 => gl_ram_ram_14(1), A2 => gl_ram_n_873, B1 => FE_OCPN151_gl_ram_ram_15_1, B2 => gl_ram_n_874, ZN => gl_ram_n_984);
  gl_ram_g8938 : AOI22D0BWP7T port map(A1 => gl_ram_ram_11(1), A2 => gl_ram_n_871, B1 => FE_OCPN72_gl_ram_ram_8_1, B2 => gl_ram_n_867, ZN => gl_ram_n_983);
  gl_ram_g8939 : AOI22D0BWP7T port map(A1 => FE_OCPN236_gl_ram_ram_82_2, A2 => gl_ram_n_868, B1 => FE_OCPN191_gl_ram_ram_83_2, B2 => gl_ram_n_871, ZN => gl_ram_n_982);
  gl_ram_g8940 : AOI22D0BWP7T port map(A1 => FE_OCPN28_gl_ram_ram_10_1, A2 => gl_ram_n_868, B1 => gl_ram_ram_9(1), B2 => gl_ram_n_869, ZN => gl_ram_n_981);
  gl_ram_g8941 : AOI22D0BWP7T port map(A1 => FE_OCPN210_gl_ram_ram_12_2, A2 => gl_ram_n_870, B1 => FE_OCPN103_gl_ram_ram_13_2, B2 => gl_ram_n_872, ZN => gl_ram_n_980);
  gl_ram_g8942 : AOI22D0BWP7T port map(A1 => FE_OCPN111_gl_ram_ram_10_2, A2 => gl_ram_n_868, B1 => gl_ram_ram_9(2), B2 => gl_ram_n_869, ZN => gl_ram_n_979);
  gl_ram_g8943 : AOI22D0BWP7T port map(A1 => gl_ram_ram_20(1), A2 => gl_ram_n_870, B1 => FE_OCPN126_gl_ram_ram_21_1, B2 => gl_ram_n_872, ZN => gl_ram_n_978);
  gl_ram_g8944 : AOI22D0BWP7T port map(A1 => gl_ram_ram_22(1), A2 => gl_ram_n_873, B1 => FE_OCPN150_gl_ram_ram_23_1, B2 => gl_ram_n_874, ZN => gl_ram_n_977);
  gl_ram_g8945 : AOI22D0BWP7T port map(A1 => FE_OCPN85_gl_ram_ram_14_2, A2 => gl_ram_n_873, B1 => FE_OCPN208_gl_ram_ram_15_2, B2 => gl_ram_n_874, ZN => gl_ram_n_976);
  gl_ram_g8946 : AOI22D0BWP7T port map(A1 => gl_ram_ram_16(1), A2 => gl_ram_n_867, B1 => gl_ram_ram_17(1), B2 => gl_ram_n_869, ZN => gl_ram_n_975);
  gl_ram_g8947 : AOI22D0BWP7T port map(A1 => gl_ram_ram_18(1), A2 => gl_ram_n_868, B1 => gl_ram_ram_19(1), B2 => gl_ram_n_871, ZN => gl_ram_n_974);
  gl_ram_g8948 : AOI22D0BWP7T port map(A1 => FE_OCPN108_gl_ram_ram_76_2, A2 => gl_ram_n_870, B1 => FE_OCPN192_gl_ram_ram_77_2, B2 => gl_ram_n_872, ZN => gl_ram_n_973);
  gl_ram_g8949 : AOI22D0BWP7T port map(A1 => gl_ram_ram_11(2), A2 => gl_ram_n_871, B1 => FE_OCPN197_gl_ram_ram_8_2, B2 => gl_ram_n_867, ZN => gl_ram_n_972);
  gl_ram_g8950 : AOI22D0BWP7T port map(A1 => FE_OCPN148_gl_ram_ram_4_1, A2 => gl_ram_n_870, B1 => gl_ram_ram_5(1), B2 => gl_ram_n_872, ZN => gl_ram_n_971);
  gl_ram_g8951 : AOI22D0BWP7T port map(A1 => gl_ram_ram_2(1), A2 => gl_ram_n_868, B1 => FE_OCPN71_gl_ram_ram_1_1, B2 => gl_ram_n_869, ZN => gl_ram_n_970);
  gl_ram_g8952 : AOI22D0BWP7T port map(A1 => FE_OCPN147_gl_ram_ram_6_1, A2 => gl_ram_n_873, B1 => gl_ram_ram_7(1), B2 => gl_ram_n_874, ZN => gl_ram_n_969);
  gl_ram_g8953 : AOI22D0BWP7T port map(A1 => gl_ram_ram_20(2), A2 => gl_ram_n_870, B1 => FE_OCPN163_gl_ram_ram_21_2, B2 => gl_ram_n_872, ZN => gl_ram_n_968);
  gl_ram_g8954 : AOI22D0BWP7T port map(A1 => FE_OCPN143_gl_ram_ram_3_1, A2 => gl_ram_n_871, B1 => FE_OCPN174_gl_ram_ram_0_1, B2 => gl_ram_n_867, ZN => gl_ram_n_967);
  gl_ram_g8955 : AOI22D0BWP7T port map(A1 => FE_OCPN214_gl_ram_ram_18_2, A2 => gl_ram_n_868, B1 => gl_ram_ram_17(2), B2 => gl_ram_n_869, ZN => gl_ram_n_966);
  gl_ram_g8956 : AOI22D0BWP7T port map(A1 => gl_ram_ram_92(0), A2 => gl_ram_n_870, B1 => gl_ram_ram_93(0), B2 => gl_ram_n_872, ZN => gl_ram_n_965);
  gl_ram_g8957 : AOI22D0BWP7T port map(A1 => gl_ram_ram_94(0), A2 => gl_ram_n_873, B1 => gl_ram_n_874, B2 => gl_ram_ram_95(0), ZN => gl_ram_n_964);
  gl_ram_g8958 : AOI22D0BWP7T port map(A1 => FE_OCPN237_gl_ram_ram_75_2, A2 => gl_ram_n_871, B1 => FE_OCPN228_gl_ram_ram_72_2, B2 => gl_ram_n_867, ZN => gl_ram_n_963);
  gl_ram_g8959 : AOI22D0BWP7T port map(A1 => FE_OCPN196_gl_ram_ram_78_2, A2 => gl_ram_n_873, B1 => FE_OCPN204_gl_ram_ram_79_2, B2 => gl_ram_n_874, ZN => gl_ram_n_962);
  gl_ram_g8960 : AOI22D0BWP7T port map(A1 => gl_ram_ram_22(2), A2 => gl_ram_n_873, B1 => FE_OCPN195_gl_ram_ram_23_2, B2 => gl_ram_n_874, ZN => gl_ram_n_961);
  gl_ram_g8961 : AOI22D0BWP7T port map(A1 => gl_ram_ram_91(0), A2 => gl_ram_n_871, B1 => gl_ram_ram_88(0), B2 => gl_ram_n_867, ZN => gl_ram_n_960);
  gl_ram_g8962 : AOI22D0BWP7T port map(A1 => gl_ram_ram_90(0), A2 => gl_ram_n_868, B1 => gl_ram_n_869, B2 => gl_ram_ram_89(0), ZN => gl_ram_n_959);
  gl_ram_g8963 : AOI22D0BWP7T port map(A1 => gl_ram_ram_19(2), A2 => gl_ram_n_871, B1 => FE_PSN355_gl_ram_ram_16_2, B2 => gl_ram_n_867, ZN => gl_ram_n_958);
  gl_ram_g8964 : AOI22D0BWP7T port map(A1 => gl_ram_ram_68(0), A2 => gl_ram_n_870, B1 => gl_ram_ram_69(0), B2 => gl_ram_n_872, ZN => gl_ram_n_957);
  gl_ram_g8965 : AOI22D0BWP7T port map(A1 => gl_ram_ram_67(0), A2 => gl_ram_n_871, B1 => gl_ram_ram_64(0), B2 => gl_ram_n_867, ZN => gl_ram_n_956);
  gl_ram_g8966 : AOI22D0BWP7T port map(A1 => gl_ram_ram_90(2), A2 => gl_ram_n_868, B1 => gl_ram_ram_89(2), B2 => gl_ram_n_869, ZN => gl_ram_n_955);
  gl_ram_g8967 : AOI22D0BWP7T port map(A1 => gl_ram_ram_74(2), A2 => gl_ram_n_868, B1 => FE_OCPN235_gl_ram_ram_73_2, B2 => gl_ram_n_869, ZN => gl_ram_n_954);
  gl_ram_g8968 : AOI22D0BWP7T port map(A1 => gl_ram_ram_4(2), A2 => gl_ram_n_870, B1 => FE_OCPN183_gl_ram_ram_5_2, B2 => gl_ram_n_872, ZN => gl_ram_n_953);
  gl_ram_g8969 : AOI22D0BWP7T port map(A1 => gl_ram_ram_70(0), A2 => gl_ram_n_873, B1 => gl_ram_ram_71(0), B2 => gl_ram_n_874, ZN => gl_ram_n_952);
  gl_ram_g8970 : AOI22D0BWP7T port map(A1 => gl_ram_ram_66(0), A2 => gl_ram_n_868, B1 => gl_ram_ram_65(0), B2 => gl_ram_n_869, ZN => gl_ram_n_951);
  gl_ram_g8971 : AOI22D0BWP7T port map(A1 => FE_OCPN194_gl_ram_ram_3_2, A2 => gl_ram_n_871, B1 => FE_OCPN221_gl_ram_ram_0_2, B2 => gl_ram_n_867, ZN => gl_ram_n_950);
  gl_ram_g8972 : AOI22D0BWP7T port map(A1 => gl_ram_ram_58(2), A2 => gl_ram_n_868, B1 => FE_OCPN169_gl_ram_ram_57_2, B2 => gl_ram_n_869, ZN => gl_ram_n_949);
  gl_ram_g8973 : AOI22D0BWP7T port map(A1 => FE_OCPN260_gl_ram_ram_2_0, A2 => gl_ram_n_868, B1 => gl_ram_ram_1(0), B2 => gl_ram_n_869, ZN => gl_ram_n_948);
  gl_ram_g8974 : AOI22D0BWP7T port map(A1 => FE_OCPN199_gl_ram_ram_2_2, A2 => gl_ram_n_868, B1 => FE_OCPN246_gl_ram_ram_1_2, B2 => gl_ram_n_869, ZN => gl_ram_n_947);
  gl_ram_g8975 : AOI22D0BWP7T port map(A1 => gl_ram_ram_84(0), A2 => gl_ram_n_870, B1 => gl_ram_ram_85(0), B2 => gl_ram_n_872, ZN => gl_ram_n_946);
  gl_ram_g8976 : AOI22D0BWP7T port map(A1 => gl_ram_ram_80(0), A2 => gl_ram_n_867, B1 => gl_ram_ram_81(0), B2 => gl_ram_n_869, ZN => gl_ram_n_945);
  gl_ram_g8977 : AOI22D0BWP7T port map(A1 => gl_ram_ram_68(2), A2 => gl_ram_n_870, B1 => FE_OCPN238_gl_ram_ram_69_2, B2 => gl_ram_n_872, ZN => gl_ram_n_944);
  gl_ram_g8978 : AOI22D0BWP7T port map(A1 => gl_ram_ram_82(0), A2 => gl_ram_n_868, B1 => gl_ram_ram_83(0), B2 => gl_ram_n_871, ZN => gl_ram_n_943);
  gl_ram_g8979 : AOI22D0BWP7T port map(A1 => gl_ram_ram_76(0), A2 => gl_ram_n_870, B1 => FE_OCPN67_gl_ram_ram_77_0, B2 => gl_ram_n_872, ZN => gl_ram_n_942);
  gl_ram_g8980 : AOI22D0BWP7T port map(A1 => FE_OCPN117_gl_ram_ram_92_1, A2 => gl_ram_n_870, B1 => gl_ram_ram_93(1), B2 => gl_ram_n_872, ZN => gl_ram_n_941);
  gl_ram_g8981 : AOI22D0BWP7T port map(A1 => gl_ram_ram_74(0), A2 => gl_ram_n_868, B1 => gl_ram_ram_73(0), B2 => gl_ram_n_869, ZN => gl_ram_n_940);
  gl_ram_g8982 : AOI22D0BWP7T port map(A1 => gl_ram_ram_52(2), A2 => gl_ram_n_870, B1 => FE_OCPN240_gl_ram_ram_53_2, B2 => gl_ram_n_872, ZN => gl_ram_n_939);
  gl_ram_g8983 : AOI22D0BWP7T port map(A1 => gl_ram_ram_94(1), A2 => gl_ram_n_873, B1 => gl_ram_ram_95(1), B2 => gl_ram_n_874, ZN => gl_ram_n_938);
  gl_ram_g8984 : AOI22D0BWP7T port map(A1 => gl_ram_ram_78(0), A2 => gl_ram_n_873, B1 => gl_ram_n_874, B2 => gl_ram_ram_79(0), ZN => gl_ram_n_937);
  gl_ram_g8985 : AOI22D0BWP7T port map(A1 => gl_ram_ram_75(0), A2 => gl_ram_n_871, B1 => gl_ram_ram_72(0), B2 => gl_ram_n_867, ZN => gl_ram_n_936);
  gl_ram_g8986 : AOI22D0BWP7T port map(A1 => FE_OCPN248_gl_ram_ram_51_2, A2 => gl_ram_n_871, B1 => FE_OCPN249_gl_ram_ram_48_2, B2 => gl_ram_n_867, ZN => gl_ram_n_935);
  gl_ram_g8987 : AOI22D0BWP7T port map(A1 => FE_OCPN145_gl_ram_ram_88_1, A2 => gl_ram_n_867, B1 => FE_OCPN140_gl_ram_ram_89_1, B2 => gl_ram_n_869, ZN => gl_ram_n_934);
  gl_ram_g8988 : AOI22D0BWP7T port map(A1 => FE_OCPN139_gl_ram_ram_90_1, A2 => gl_ram_n_868, B1 => FE_OCPN119_gl_ram_ram_91_1, B2 => gl_ram_n_871, ZN => gl_ram_n_933);
  gl_ram_g8989 : AOI22D0BWP7T port map(A1 => FE_OCPN42_gl_ram_ram_60_0, A2 => gl_ram_n_870, B1 => gl_ram_ram_61(0), B2 => gl_ram_n_872, ZN => gl_ram_n_932);
  gl_ram_g8990 : AOI22D0BWP7T port map(A1 => gl_ram_ram_59(0), A2 => gl_ram_n_871, B1 => FE_OCPN43_gl_ram_ram_56_0, B2 => gl_ram_n_867, ZN => gl_ram_n_931);
  gl_ram_g8991 : AOI22D0BWP7T port map(A1 => gl_ram_ram_62(0), A2 => gl_ram_n_873, B1 => FE_OCPN267_gl_ram_ram_63_0, B2 => gl_ram_n_874, ZN => gl_ram_n_930);
  gl_ram_g8992 : AOI22D0BWP7T port map(A1 => gl_ram_ram_66(2), A2 => gl_ram_n_868, B1 => FE_OCPN198_gl_ram_ram_65_2, B2 => gl_ram_n_869, ZN => gl_ram_n_929);
  gl_ram_g8993 : AOI22D0BWP7T port map(A1 => gl_ram_ram_58(0), A2 => gl_ram_n_868, B1 => gl_ram_n_869, B2 => gl_ram_ram_57(0), ZN => gl_ram_n_928);
  gl_ram_g8994 : AOI22D0BWP7T port map(A1 => gl_ram_ram_54(2), A2 => gl_ram_n_873, B1 => FE_OCPN61_gl_ram_ram_55_2, B2 => gl_ram_n_874, ZN => gl_ram_n_927);
  gl_ram_g8995 : AOI22D0BWP7T port map(A1 => gl_ram_ram_68(1), A2 => gl_ram_n_870, B1 => gl_ram_ram_69(1), B2 => gl_ram_n_872, ZN => gl_ram_n_926);
  gl_ram_g8996 : AOI22D0BWP7T port map(A1 => gl_ram_ram_36(0), A2 => gl_ram_n_870, B1 => FE_OCPN175_gl_ram_ram_37_0, B2 => gl_ram_n_872, ZN => gl_ram_n_925);
  gl_ram_g8997 : AOI22D0BWP7T port map(A1 => gl_ram_ram_38(0), A2 => gl_ram_n_873, B1 => gl_ram_ram_39(0), B2 => gl_ram_n_874, ZN => gl_ram_n_924);
  gl_ram_g8998 : AOI22D0BWP7T port map(A1 => gl_ram_ram_66(1), A2 => gl_ram_n_868, B1 => gl_ram_ram_65(1), B2 => gl_ram_n_869, ZN => gl_ram_n_923);
  gl_ram_g8999 : AOI22D0BWP7T port map(A1 => gl_ram_ram_35(0), A2 => gl_ram_n_871, B1 => gl_ram_ram_32(0), B2 => gl_ram_n_867, ZN => gl_ram_n_922);
  gl_ram_g9000 : AOI22D0BWP7T port map(A1 => FE_OCPN231_gl_ram_ram_50_2, A2 => gl_ram_n_868, B1 => gl_ram_ram_49(2), B2 => gl_ram_n_869, ZN => gl_ram_n_921);
  gl_ram_g9001 : AOI22D0BWP7T port map(A1 => gl_ram_ram_34(0), A2 => gl_ram_n_868, B1 => gl_ram_ram_33(0), B2 => gl_ram_n_869, ZN => gl_ram_n_920);
  gl_ram_g9002 : AOI22D0BWP7T port map(A1 => gl_ram_ram_70(1), A2 => gl_ram_n_873, B1 => FE_OCPN116_gl_ram_ram_71_1, B2 => gl_ram_n_874, ZN => gl_ram_n_919);
  gl_ram_g9003 : AOI22D0BWP7T port map(A1 => gl_ram_ram_70(2), A2 => gl_ram_n_873, B1 => FE_OCPN218_gl_ram_ram_71_2, B2 => gl_ram_n_874, ZN => gl_ram_n_918);
  gl_ram_g9004 : AOI22D0BWP7T port map(A1 => FE_OCPN243_gl_ram_ram_28_0, A2 => gl_ram_n_870, B1 => FE_OCPN66_gl_ram_ram_29_0, B2 => gl_ram_n_872, ZN => gl_ram_n_917);
  gl_ram_g9005 : AOI22D0BWP7T port map(A1 => FE_OCPN125_gl_ram_ram_67_1, A2 => gl_ram_n_871, B1 => gl_ram_ram_64(1), B2 => gl_ram_n_867, ZN => gl_ram_n_916);
  gl_ram_g9006 : AOI22D0BWP7T port map(A1 => FE_OCPN264_gl_ram_ram_30_0, A2 => gl_ram_n_873, B1 => FE_OCPN63_gl_ram_ram_31_0, B2 => gl_ram_n_874, ZN => gl_ram_n_915);
  gl_ram_g9007 : AOI22D0BWP7T port map(A1 => FE_OCPN193_gl_ram_ram_92_2, A2 => gl_ram_n_870, B1 => gl_ram_ram_93(2), B2 => gl_ram_n_872, ZN => gl_ram_n_914);
  gl_ram_g9008 : AOI22D0BWP7T port map(A1 => gl_ram_ram_27(0), A2 => gl_ram_n_871, B1 => FE_OCPN89_gl_ram_ram_24_0, B2 => gl_ram_n_867, ZN => gl_ram_n_913);
  gl_ram_g9009 : AOI22D0BWP7T port map(A1 => FE_OCPN217_gl_ram_ram_67_2, A2 => gl_ram_n_871, B1 => gl_ram_ram_64(2), B2 => gl_ram_n_867, ZN => gl_ram_n_912);
  gl_ram_g9010 : AOI22D0BWP7T port map(A1 => gl_ram_ram_26(0), A2 => gl_ram_n_868, B1 => gl_ram_n_869, B2 => gl_ram_ram_25(0), ZN => gl_ram_n_911);
  gl_ram_g9011 : AOI22D0BWP7T port map(A1 => gl_ram_ram_91(2), A2 => gl_ram_n_871, B1 => gl_ram_ram_88(2), B2 => gl_ram_n_867, ZN => gl_ram_n_910);
  gl_ram_g9012 : AOI22D0BWP7T port map(A1 => gl_ram_ram_12(0), A2 => gl_ram_n_870, B1 => FE_OCPN186_gl_ram_ram_13_0, B2 => gl_ram_n_872, ZN => gl_ram_n_909);
  gl_ram_g9013 : AOI22D0BWP7T port map(A1 => FE_OCPN203_gl_ram_ram_44_2, A2 => gl_ram_n_870, B1 => gl_ram_n_872, B2 => gl_ram_ram_45(2), ZN => gl_ram_n_908);
  gl_ram_g9014 : AOI22D0BWP7T port map(A1 => gl_ram_ram_14(0), A2 => gl_ram_n_873, B1 => FE_OCPN255_gl_ram_ram_15_0, B2 => gl_ram_n_874, ZN => gl_ram_n_907);
  gl_ram_g9015 : AOI22D0BWP7T port map(A1 => gl_ram_ram_11(0), A2 => gl_ram_n_871, B1 => gl_ram_ram_8(0), B2 => gl_ram_n_867, ZN => gl_ram_n_906);
  gl_ram_g9016 : AOI22D0BWP7T port map(A1 => FE_OCPN268_gl_ram_ram_10_0, A2 => gl_ram_n_868, B1 => FE_OCPN259_gl_ram_ram_9_0, B2 => gl_ram_n_869, ZN => gl_ram_n_905);
  gl_ram_g9017 : AOI22D0BWP7T port map(A1 => FE_OCPN189_gl_ram_ram_52_0, A2 => gl_ram_n_870, B1 => gl_ram_ram_53(0), B2 => gl_ram_n_872, ZN => gl_ram_n_904);
  gl_ram_g9018 : AOI22D0BWP7T port map(A1 => gl_ram_ram_50(0), A2 => gl_ram_n_868, B1 => FE_OCPN262_gl_ram_ram_49_0, B2 => gl_ram_n_869, ZN => gl_ram_n_903);
  gl_ram_g9019 : AO22D0BWP7T port map(A1 => gl_ram_ram_98(1), A2 => gl_ram_n_868, B1 => gl_ram_n_871, B2 => gl_ram_ram_99(1), Z => gl_ram_n_902);
  gl_ram_g9020 : AOI22D0BWP7T port map(A1 => gl_ram_ram_84(1), A2 => gl_ram_n_870, B1 => FE_OCPN123_gl_ram_ram_85_1, B2 => gl_ram_n_872, ZN => gl_ram_n_901);
  gl_ram_g9021 : AOI22D0BWP7T port map(A1 => FE_OCPN265_gl_ram_ram_54_0, A2 => gl_ram_n_873, B1 => FE_OCPN266_gl_ram_ram_55_0, B2 => gl_ram_n_874, ZN => gl_ram_n_900);
  gl_ram_g9022 : AOI22D0BWP7T port map(A1 => gl_ram_ram_51(0), A2 => gl_ram_n_871, B1 => FE_OCPN38_gl_ram_ram_48_0, B2 => gl_ram_n_867, ZN => gl_ram_n_899);
  gl_ram_g9023 : AOI22D0BWP7T port map(A1 => gl_ram_ram_43(2), A2 => gl_ram_n_871, B1 => FE_OCPN271_gl_ram_ram_40_2, B2 => gl_ram_n_867, ZN => gl_ram_n_898);
  gl_ram_g9024 : AOI22D0BWP7T port map(A1 => gl_ram_ram_83(1), A2 => gl_ram_n_871, B1 => FE_OCPN130_gl_ram_ram_80_1, B2 => gl_ram_n_867, ZN => gl_ram_n_897);
  gl_ram_g9025 : AOI22D0BWP7T port map(A1 => FE_OCPN226_gl_ram_ram_46_2, A2 => gl_ram_n_873, B1 => gl_ram_n_874, B2 => FE_OCPN200_gl_ram_ram_47_2, ZN => gl_ram_n_896);
  gl_ram_g9026 : AOI22D0BWP7T port map(A1 => gl_ram_ram_44(0), A2 => gl_ram_n_870, B1 => gl_ram_ram_45(0), B2 => gl_ram_n_872, ZN => gl_ram_n_895);
  gl_ram_g9027 : AOI22D0BWP7T port map(A1 => FE_OCPN272_gl_ram_ram_43_0, A2 => gl_ram_n_871, B1 => FE_OCPN170_gl_ram_ram_40_0, B2 => gl_ram_n_867, ZN => gl_ram_n_894);
  gl_ram_g9028 : AOI22D0BWP7T port map(A1 => gl_ram_ram_82(1), A2 => gl_ram_n_868, B1 => FE_OCPN127_gl_ram_ram_81_1, B2 => gl_ram_n_869, ZN => gl_ram_n_893);
  gl_ram_g9029 : AOI22D0BWP7T port map(A1 => gl_ram_ram_46(0), A2 => gl_ram_n_873, B1 => gl_ram_ram_47(0), B2 => gl_ram_n_874, ZN => gl_ram_n_892);
  gl_ram_g9030 : AOI22D0BWP7T port map(A1 => gl_ram_ram_42(2), A2 => gl_ram_n_868, B1 => FE_OCPN247_gl_ram_ram_41_2, B2 => gl_ram_n_869, ZN => gl_ram_n_891);
  gl_ram_g9031 : AOI22D0BWP7T port map(A1 => FE_OCPN257_gl_ram_ram_42_0, A2 => gl_ram_n_868, B1 => FE_OCPN46_gl_ram_ram_41_0, B2 => gl_ram_n_869, ZN => gl_ram_n_890);
  gl_ram_g9032 : AOI22D0BWP7T port map(A1 => gl_ram_ram_20(0), A2 => gl_ram_n_870, B1 => FE_OCPN74_gl_ram_ram_21_0, B2 => gl_ram_n_872, ZN => gl_ram_n_889);
  gl_ram_g9033 : AOI22D0BWP7T port map(A1 => FE_OCPN133_gl_ram_ram_76_1, A2 => gl_ram_n_870, B1 => FE_OCPN110_gl_ram_ram_77_1, B2 => gl_ram_n_872, ZN => gl_ram_n_888);
  gl_ram_g9034 : AOI22D0BWP7T port map(A1 => gl_ram_ram_19(0), A2 => gl_ram_n_871, B1 => gl_ram_ram_16(0), B2 => gl_ram_n_867, ZN => gl_ram_n_887);
  gl_ram_g9035 : AOI22D0BWP7T port map(A1 => FE_OCPN65_gl_ram_ram_74_1, A2 => gl_ram_n_868, B1 => FE_OCPN70_gl_ram_ram_73_1, B2 => gl_ram_n_869, ZN => gl_ram_n_886);
  gl_ram_g9036 : AOI22D0BWP7T port map(A1 => gl_ram_ram_22(0), A2 => gl_ram_n_873, B1 => gl_ram_n_874, B2 => gl_ram_ram_23(0), ZN => gl_ram_n_885);
  gl_ram_g9037 : AOI22D0BWP7T port map(A1 => gl_ram_ram_18(0), A2 => gl_ram_n_868, B1 => gl_ram_ram_17(0), B2 => gl_ram_n_869, ZN => gl_ram_n_884);
  gl_ram_g9038 : AOI22D0BWP7T port map(A1 => FE_OCPN107_gl_ram_ram_78_1, A2 => gl_ram_n_873, B1 => FE_OCPN102_gl_ram_ram_79_1, B2 => gl_ram_n_874, ZN => gl_ram_n_883);
  gl_ram_g9039 : AOI22D0BWP7T port map(A1 => FE_OCPN263_gl_ram_ram_4_0, A2 => gl_ram_n_870, B1 => FE_OCPN245_gl_ram_ram_5_0, B2 => gl_ram_n_872, ZN => gl_ram_n_882);
  gl_ram_g9040 : AOI22D0BWP7T port map(A1 => gl_ram_ram_3(0), A2 => gl_ram_n_871, B1 => gl_ram_ram_0(0), B2 => gl_ram_n_867, ZN => gl_ram_n_881);
  gl_ram_g9041 : AOI22D0BWP7T port map(A1 => gl_ram_ram_60(2), A2 => gl_ram_n_870, B1 => gl_ram_ram_61(2), B2 => gl_ram_n_872, ZN => gl_ram_n_880);
  gl_ram_g9042 : AOI22D0BWP7T port map(A1 => gl_ram_ram_75(1), A2 => gl_ram_n_871, B1 => gl_ram_ram_72(1), B2 => gl_ram_n_867, ZN => gl_ram_n_879);
  gl_ram_g9043 : AOI22D0BWP7T port map(A1 => gl_ram_ram_6(0), A2 => gl_ram_n_873, B1 => gl_ram_ram_7(0), B2 => gl_ram_n_874, ZN => gl_ram_n_878);
  gl_ram_g9044 : AOI22D0BWP7T port map(A1 => FE_OCPN180_gl_ram_ram_6_2, A2 => gl_ram_n_873, B1 => FE_OCPN173_gl_ram_ram_7_2, B2 => gl_ram_n_874, ZN => gl_ram_n_877);
  gl_ram_g9045 : FA1D0BWP7T port map(A => gl_ram_n_858, B => gl_sig_y(2), CI => gl_ram_n_859, CO => gl_ram_n_875, S => gl_ram_n_876);
  gl_ram_g9047 : AN2D1BWP7T port map(A1 => gl_ram_n_863, A2 => gl_sig_x(0), Z => gl_ram_n_874);
  gl_ram_g9048 : NR2XD1BWP7T port map(A1 => gl_ram_n_862, A2 => gl_sig_x(0), ZN => gl_ram_n_873);
  gl_ram_g9049 : INR2XD2BWP7T port map(A1 => gl_sig_x(0), B1 => gl_ram_n_861, ZN => gl_ram_n_872);
  gl_ram_g9050 : CKAN2D2BWP7T port map(A1 => gl_ram_n_864, A2 => gl_sig_x(0), Z => gl_ram_n_871);
  gl_ram_g9051 : NR2D2P5BWP7T port map(A1 => gl_ram_n_861, A2 => gl_sig_x(0), ZN => gl_ram_n_870);
  gl_ram_g9052 : CKAN2D2BWP7T port map(A1 => gl_ram_n_866, A2 => gl_sig_x(0), Z => gl_ram_n_869);
  gl_ram_g9053 : INR2XD2BWP7T port map(A1 => gl_ram_n_864, B1 => gl_sig_x(0), ZN => gl_ram_n_868);
  gl_ram_g9054 : NR2D2P5BWP7T port map(A1 => gl_ram_n_865, A2 => gl_sig_x(0), ZN => gl_ram_n_867);
  gl_ram_g9055 : INVD0BWP7T port map(I => gl_ram_n_865, ZN => gl_ram_n_866);
  gl_ram_g9056 : IND2D1BWP7T port map(A1 => gl_ram_n_860, B1 => gl_ram_n_842, ZN => gl_ram_n_865);
  gl_ram_g9057 : NR2D1BWP7T port map(A1 => gl_ram_n_860, A2 => gl_ram_n_842, ZN => gl_ram_n_864);
  gl_ram_g9058 : INVD1BWP7T port map(I => gl_ram_n_862, ZN => gl_ram_n_863);
  gl_ram_g9059 : IND2D1BWP7T port map(A1 => gl_ram_n_842, B1 => gl_ram_n_860, ZN => gl_ram_n_862);
  gl_ram_g9060 : ND2D1BWP7T port map(A1 => gl_ram_n_860, A2 => gl_ram_n_842, ZN => gl_ram_n_861);
  gl_ram_g9061 : FA1D0BWP7T port map(A => gl_sig_y(1), B => gl_sig_x(2), CI => gl_ram_n_824, CO => gl_ram_n_859, S => gl_ram_n_860);
  gl_ram_g9062 : NR2D0BWP7T port map(A1 => gl_ram_n_854, A2 => gl_ram_n_844, ZN => gl_ram_n_1110);
  gl_ram_g9063 : NR2D0BWP7T port map(A1 => gl_ram_n_854, A2 => gl_ram_n_843, ZN => gl_ram_n_1116);
  gl_ram_g9064 : NR2D0BWP7T port map(A1 => gl_ram_n_854, A2 => gl_ram_n_845, ZN => gl_ram_n_1114);
  gl_ram_g9065 : NR2D0BWP7T port map(A1 => gl_ram_n_854, A2 => gl_ram_n_833, ZN => gl_ram_n_1112);
  gl_ram_g9066 : HA1D0BWP7T port map(A => gl_sig_x(3), B => gl_sig_y(0), CO => gl_ram_n_857, S => gl_ram_n_858);
  gl_ram_g9067 : HA1D0BWP7T port map(A => gl_sig_y(3), B => gl_sig_y(1), CO => gl_ram_n_855, S => gl_ram_n_856);
  gl_ram_g9068 : NR2D0BWP7T port map(A1 => gl_ram_n_853, A2 => gl_ram_n_847, ZN => gl_ram_n_1262);
  gl_ram_g9069 : NR2D0BWP7T port map(A1 => gl_ram_n_851, A2 => gl_ram_n_834, ZN => gl_ram_n_1296);
  gl_ram_g9070 : NR2D0BWP7T port map(A1 => gl_ram_n_840, A2 => gl_ram_n_834, ZN => gl_ram_n_1280);
  gl_ram_g9071 : NR2D0BWP7T port map(A1 => gl_ram_n_853, A2 => gl_ram_n_834, ZN => gl_ram_n_1264);
  gl_ram_g9072 : NR2D0BWP7T port map(A1 => gl_ram_n_849, A2 => gl_ram_n_834, ZN => gl_ram_n_1232);
  gl_ram_g9073 : NR2D0BWP7T port map(A1 => gl_ram_n_850, A2 => gl_ram_n_835, ZN => gl_ram_n_1186);
  gl_ram_g9074 : NR2D0BWP7T port map(A1 => gl_ram_n_850, A2 => gl_ram_n_846, ZN => gl_ram_n_1188);
  gl_ram_g9075 : NR2D0BWP7T port map(A1 => gl_ram_n_848, A2 => gl_ram_n_846, ZN => gl_ram_n_1124);
  gl_ram_g9076 : NR2D0BWP7T port map(A1 => gl_ram_n_848, A2 => gl_ram_n_835, ZN => gl_ram_n_1122);
  gl_ram_g9077 : NR2D0BWP7T port map(A1 => gl_ram_n_838, A2 => gl_ram_n_834, ZN => gl_ram_n_1168);
  gl_ram_g9078 : NR2D0BWP7T port map(A1 => gl_ram_n_851, A2 => gl_ram_n_833, ZN => gl_ram_n_1304);
  gl_ram_g9079 : NR2D0BWP7T port map(A1 => gl_ram_n_851, A2 => gl_ram_n_844, ZN => gl_ram_n_1302);
  gl_ram_g9080 : NR2D0BWP7T port map(A1 => gl_ram_n_853, A2 => gl_ram_n_833, ZN => gl_ram_n_1272);
  gl_ram_g9081 : NR2D0BWP7T port map(A1 => gl_ram_n_849, A2 => gl_ram_n_833, ZN => gl_ram_n_1240);
  gl_ram_g9082 : NR2D0BWP7T port map(A1 => gl_ram_n_850, A2 => gl_ram_n_845, ZN => gl_ram_n_1194);
  gl_ram_g9083 : NR2D0BWP7T port map(A1 => gl_ram_n_838, A2 => gl_ram_n_833, ZN => gl_ram_n_1176);
  gl_ram_g9084 : NR2D0BWP7T port map(A1 => gl_ram_n_838, A2 => gl_ram_n_844, ZN => gl_ram_n_1174);
  gl_ram_g9085 : NR2D0BWP7T port map(A1 => gl_ram_n_848, A2 => gl_ram_n_845, ZN => gl_ram_n_1130);
  gl_ram_g9086 : NR2D0BWP7T port map(A1 => gl_ram_n_853, A2 => gl_ram_n_844, ZN => gl_ram_n_1270);
  gl_ram_g9087 : NR2D0BWP7T port map(A1 => gl_ram_n_840, A2 => gl_ram_n_833, ZN => gl_ram_n_1288);
  gl_ram_g9088 : NR2D0BWP7T port map(A1 => gl_ram_n_840, A2 => gl_ram_n_844, ZN => gl_ram_n_1286);
  gl_ram_g9089 : NR2D0BWP7T port map(A1 => gl_ram_n_849, A2 => gl_ram_n_844, ZN => gl_ram_n_1238);
  gl_ram_g9090 : NR2D0BWP7T port map(A1 => gl_ram_n_838, A2 => gl_ram_n_835, ZN => gl_ram_n_1170);
  gl_ram_g9091 : NR2D0BWP7T port map(A1 => gl_ram_n_851, A2 => gl_ram_n_843, ZN => gl_ram_n_1308);
  gl_ram_g9092 : NR2D0BWP7T port map(A1 => gl_ram_n_851, A2 => gl_ram_n_845, ZN => gl_ram_n_1306);
  gl_ram_g9093 : NR2D0BWP7T port map(A1 => gl_ram_n_851, A2 => gl_ram_n_835, ZN => gl_ram_n_1298);
  gl_ram_g9094 : NR2D0BWP7T port map(A1 => gl_ram_n_840, A2 => gl_ram_n_843, ZN => gl_ram_n_1292);
  gl_ram_g9095 : NR2D0BWP7T port map(A1 => gl_ram_n_840, A2 => gl_ram_n_845, ZN => gl_ram_n_1290);
  gl_ram_g9096 : NR2D0BWP7T port map(A1 => gl_ram_n_840, A2 => gl_ram_n_846, ZN => gl_ram_n_1284);
  gl_ram_g9097 : NR2D0BWP7T port map(A1 => gl_ram_n_853, A2 => gl_ram_n_843, ZN => gl_ram_n_1276);
  gl_ram_g9098 : NR2D0BWP7T port map(A1 => gl_ram_n_853, A2 => gl_ram_n_845, ZN => gl_ram_n_1274);
  gl_ram_g9099 : NR2D0BWP7T port map(A1 => gl_ram_n_853, A2 => gl_ram_n_846, ZN => gl_ram_n_1268);
  gl_ram_g9100 : NR2D0BWP7T port map(A1 => gl_ram_n_849, A2 => gl_ram_n_843, ZN => gl_ram_n_1244);
  gl_ram_g9101 : NR2D0BWP7T port map(A1 => gl_ram_n_849, A2 => gl_ram_n_845, ZN => gl_ram_n_1242);
  gl_ram_g9102 : NR2D0BWP7T port map(A1 => gl_ram_n_849, A2 => gl_ram_n_846, ZN => gl_ram_n_1236);
  gl_ram_g9103 : NR2D0BWP7T port map(A1 => gl_ram_n_849, A2 => gl_ram_n_847, ZN => gl_ram_n_1230);
  gl_ram_g9104 : NR2D0BWP7T port map(A1 => gl_ram_n_850, A2 => gl_ram_n_847, ZN => gl_ram_n_1182);
  gl_ram_g9105 : NR2D0BWP7T port map(A1 => gl_ram_n_850, A2 => gl_ram_n_833, ZN => gl_ram_n_1192);
  gl_ram_g9106 : NR2D0BWP7T port map(A1 => gl_ram_n_838, A2 => gl_ram_n_847, ZN => gl_ram_n_1166);
  gl_ram_g9107 : NR2D0BWP7T port map(A1 => gl_ram_n_848, A2 => gl_ram_n_843, ZN => gl_ram_n_1132);
  gl_ram_g9108 : NR2D0BWP7T port map(A1 => gl_ram_n_848, A2 => gl_ram_n_833, ZN => gl_ram_n_1128);
  gl_ram_g9109 : NR2D0BWP7T port map(A1 => gl_ram_n_851, A2 => gl_ram_n_847, ZN => gl_ram_n_1294);
  gl_ram_g9110 : NR2D0BWP7T port map(A1 => gl_ram_n_848, A2 => gl_ram_n_844, ZN => gl_ram_n_1126);
  gl_ram_g9111 : NR2D0BWP7T port map(A1 => gl_ram_n_850, A2 => gl_ram_n_843, ZN => gl_ram_n_1196);
  gl_ram_g9112 : NR2D0BWP7T port map(A1 => gl_ram_n_848, A2 => gl_ram_n_847, ZN => gl_ram_n_1118);
  gl_ram_g9113 : NR2D0BWP7T port map(A1 => gl_ram_n_849, A2 => gl_ram_n_835, ZN => gl_ram_n_1234);
  gl_ram_g9114 : NR2D0BWP7T port map(A1 => gl_ram_n_848, A2 => gl_ram_n_834, ZN => gl_ram_n_1120);
  gl_ram_g9115 : NR2D0BWP7T port map(A1 => gl_ram_n_838, A2 => gl_ram_n_845, ZN => gl_ram_n_1178);
  gl_ram_g9116 : AOI21D2BWP7T port map(A1 => FE_PHN292_gl_ram_n_819, A2 => FE_PHN291_gl_ram_n_1310, B => gl_ram_n_1320, ZN => gl_ram_n_1111);
  gl_ram_g9117 : NR2D0BWP7T port map(A1 => gl_ram_n_850, A2 => gl_ram_n_844, ZN => gl_ram_n_1190);
  gl_ram_g9118 : NR2D0BWP7T port map(A1 => gl_ram_n_840, A2 => gl_ram_n_835, ZN => gl_ram_n_1282);
  gl_ram_g9119 : NR2D0BWP7T port map(A1 => gl_ram_n_838, A2 => gl_ram_n_843, ZN => gl_ram_n_1180);
  gl_ram_g9120 : NR2D0BWP7T port map(A1 => gl_ram_n_853, A2 => gl_ram_n_835, ZN => gl_ram_n_1266);
  gl_ram_g9121 : NR2D0BWP7T port map(A1 => gl_ram_n_840, A2 => gl_ram_n_847, ZN => gl_ram_n_1278);
  gl_ram_g9122 : NR2D0BWP7T port map(A1 => gl_ram_n_838, A2 => gl_ram_n_846, ZN => gl_ram_n_1172);
  gl_ram_g9123 : NR2D0BWP7T port map(A1 => gl_ram_n_851, A2 => gl_ram_n_846, ZN => gl_ram_n_1300);
  gl_ram_g9124 : NR2D0BWP7T port map(A1 => gl_ram_n_852, A2 => gl_ram_n_846, ZN => gl_ram_n_1252);
  gl_ram_g9125 : NR2D0BWP7T port map(A1 => gl_ram_n_852, A2 => gl_ram_n_834, ZN => gl_ram_n_1248);
  gl_ram_g9126 : NR2D0BWP7T port map(A1 => gl_ram_n_841, A2 => gl_ram_n_846, ZN => gl_ram_n_1220);
  gl_ram_g9127 : NR2D0BWP7T port map(A1 => gl_ram_n_836, A2 => gl_ram_n_834, ZN => gl_ram_n_1200);
  gl_ram_g9128 : NR2D0BWP7T port map(A1 => gl_ram_n_837, A2 => gl_ram_n_835, ZN => gl_ram_n_1154);
  gl_ram_g9129 : NR2D0BWP7T port map(A1 => gl_ram_n_837, A2 => gl_ram_n_834, ZN => gl_ram_n_1152);
  gl_ram_g9130 : NR2D0BWP7T port map(A1 => gl_ram_n_839, A2 => gl_ram_n_835, ZN => gl_ram_n_1138);
  gl_ram_g9131 : NR2D0BWP7T port map(A1 => gl_ram_n_841, A2 => gl_ram_n_835, ZN => gl_ram_n_1218);
  gl_ram_g9132 : NR2D0BWP7T port map(A1 => gl_ram_n_836, A2 => gl_ram_n_846, ZN => gl_ram_n_1204);
  gl_ram_g9133 : NR2D0BWP7T port map(A1 => gl_ram_n_837, A2 => gl_ram_n_846, ZN => gl_ram_n_1156);
  gl_ram_g9134 : NR2D0BWP7T port map(A1 => gl_ram_n_839, A2 => gl_ram_n_834, ZN => gl_ram_n_1136);
  gl_ram_g9135 : NR2D0BWP7T port map(A1 => gl_ram_n_839, A2 => gl_ram_n_846, ZN => gl_ram_n_1140);
  gl_ram_g9136 : NR2D0BWP7T port map(A1 => gl_ram_n_841, A2 => gl_ram_n_834, ZN => gl_ram_n_1216);
  gl_ram_g9137 : NR2D0BWP7T port map(A1 => gl_ram_n_852, A2 => gl_ram_n_835, ZN => gl_ram_n_1250);
  gl_ram_g9138 : NR2D0BWP7T port map(A1 => gl_ram_n_836, A2 => gl_ram_n_835, ZN => gl_ram_n_1202);
  gl_ram_g9139 : NR2D0BWP7T port map(A1 => gl_ram_n_837, A2 => gl_ram_n_845, ZN => gl_ram_n_1162);
  gl_ram_g9140 : NR2D0BWP7T port map(A1 => gl_ram_n_852, A2 => gl_ram_n_845, ZN => gl_ram_n_1258);
  gl_ram_g9141 : NR2D0BWP7T port map(A1 => gl_ram_n_841, A2 => gl_ram_n_845, ZN => gl_ram_n_1226);
  gl_ram_g9142 : NR2D0BWP7T port map(A1 => gl_ram_n_836, A2 => gl_ram_n_845, ZN => gl_ram_n_1210);
  gl_ram_g9143 : NR2D0BWP7T port map(A1 => gl_ram_n_839, A2 => gl_ram_n_844, ZN => gl_ram_n_1142);
  gl_ram_g9144 : NR2D0BWP7T port map(A1 => gl_ram_n_837, A2 => gl_ram_n_833, ZN => gl_ram_n_1160);
  gl_ram_g9145 : NR2D0BWP7T port map(A1 => gl_ram_n_839, A2 => gl_ram_n_845, ZN => gl_ram_n_1146);
  gl_ram_g9146 : NR2D0BWP7T port map(A1 => gl_ram_n_852, A2 => gl_ram_n_844, ZN => gl_ram_n_1254);
  gl_ram_g9147 : NR2D0BWP7T port map(A1 => gl_ram_n_836, A2 => gl_ram_n_833, ZN => gl_ram_n_1208);
  gl_ram_g9148 : NR2D0BWP7T port map(A1 => gl_ram_n_841, A2 => gl_ram_n_833, ZN => gl_ram_n_1224);
  gl_ram_g9149 : NR2D0BWP7T port map(A1 => gl_ram_n_836, A2 => gl_ram_n_844, ZN => gl_ram_n_1206);
  gl_ram_g9150 : NR2D0BWP7T port map(A1 => gl_ram_n_837, A2 => gl_ram_n_844, ZN => gl_ram_n_1158);
  gl_ram_g9151 : NR2D0BWP7T port map(A1 => gl_ram_n_841, A2 => gl_ram_n_844, ZN => gl_ram_n_1222);
  gl_ram_g9152 : NR2D0BWP7T port map(A1 => gl_ram_n_852, A2 => gl_ram_n_833, ZN => gl_ram_n_1256);
  gl_ram_g9153 : NR2D0BWP7T port map(A1 => gl_ram_n_839, A2 => gl_ram_n_833, ZN => gl_ram_n_1144);
  gl_ram_g9154 : NR2D0BWP7T port map(A1 => gl_ram_n_852, A2 => gl_ram_n_847, ZN => gl_ram_n_1246);
  gl_ram_g9155 : NR2D0BWP7T port map(A1 => gl_ram_n_841, A2 => gl_ram_n_847, ZN => gl_ram_n_1214);
  gl_ram_g9156 : NR2D0BWP7T port map(A1 => gl_ram_n_839, A2 => gl_ram_n_843, ZN => gl_ram_n_1148);
  gl_ram_g9157 : NR2D0BWP7T port map(A1 => gl_ram_n_837, A2 => gl_ram_n_847, ZN => gl_ram_n_1150);
  gl_ram_g9158 : NR2D0BWP7T port map(A1 => gl_ram_n_836, A2 => gl_ram_n_847, ZN => gl_ram_n_1198);
  gl_ram_g9159 : NR2D0BWP7T port map(A1 => gl_ram_n_839, A2 => gl_ram_n_847, ZN => gl_ram_n_1134);
  gl_ram_g9160 : NR2D0BWP7T port map(A1 => gl_ram_n_837, A2 => gl_ram_n_843, ZN => gl_ram_n_1164);
  gl_ram_g9161 : NR2D0BWP7T port map(A1 => gl_ram_n_836, A2 => gl_ram_n_843, ZN => gl_ram_n_1212);
  gl_ram_g9162 : NR2D0BWP7T port map(A1 => gl_ram_n_841, A2 => gl_ram_n_843, ZN => gl_ram_n_1228);
  gl_ram_g9163 : NR2D0BWP7T port map(A1 => gl_ram_n_852, A2 => gl_ram_n_843, ZN => gl_ram_n_1260);
  gl_ram_g9164 : NR2D0BWP7T port map(A1 => gl_ram_n_850, A2 => gl_ram_n_834, ZN => gl_ram_n_1184);
  gl_ram_g9165 : ND3D0BWP7T port map(A1 => gl_ram_n_821, A2 => gl_ram_ram_position(6), A3 => gl_ram_ram_position(5), ZN => gl_ram_n_854);
  gl_ram_g9166 : ND2D0BWP7T port map(A1 => gl_ram_n_829, A2 => gl_ram_n_822, ZN => gl_ram_n_853);
  gl_ram_g9167 : IND2D0BWP7T port map(A1 => gl_ram_n_828, B1 => gl_ram_n_822, ZN => gl_ram_n_852);
  gl_ram_g9168 : ND2D0BWP7T port map(A1 => gl_ram_n_821, A2 => gl_ram_n_822, ZN => gl_ram_n_851);
  gl_ram_g9169 : IND2D0BWP7T port map(A1 => gl_ram_n_828, B1 => gl_ram_n_820, ZN => gl_ram_n_850);
  gl_ram_g9170 : ND2D0BWP7T port map(A1 => gl_ram_n_820, A2 => gl_ram_n_821, ZN => gl_ram_n_849);
  gl_ram_g9171 : IND2D0BWP7T port map(A1 => gl_ram_n_828, B1 => gl_ram_n_827, ZN => gl_ram_n_848);
  gl_ram_g9172 : IND2D1BWP7T port map(A1 => gl_ram_n_832, B1 => gl_ram_ram_position(1), ZN => gl_ram_n_847);
  gl_ram_g9173 : IND2D1BWP7T port map(A1 => gl_ram_ram_position(1), B1 => gl_ram_n_830, ZN => gl_ram_n_846);
  gl_ram_g9174 : IND2D1BWP7T port map(A1 => gl_ram_ram_position(1), B1 => gl_ram_n_826, ZN => gl_ram_n_845);
  gl_ram_g9175 : CKND2D1BWP7T port map(A1 => gl_ram_n_826, A2 => gl_ram_ram_position(1), ZN => gl_ram_n_844);
  gl_ram_g9176 : IND2D1BWP7T port map(A1 => gl_ram_ram_position(1), B1 => gl_ram_n_831, ZN => gl_ram_n_843);
  gl_ram_g9177 : INR3D0BWP7T port map(A1 => FE_PHN294_gl_ram_n_1311, B1 => FE_PHN314_sig_logic_x_3, B2 => FE_PHN286_sig_logic_x_2, ZN => gl_ram_n_1320);
  gl_ram_g9178 : OAI21D0BWP7T port map(A1 => gl_sig_y(0), A2 => gl_sig_x(1), B => gl_ram_n_823, ZN => gl_ram_n_842);
  gl_ram_g9179 : ND2D0BWP7T port map(A1 => gl_ram_n_820, A2 => gl_ram_n_825, ZN => gl_ram_n_841);
  gl_ram_g9180 : ND2D0BWP7T port map(A1 => gl_ram_n_825, A2 => gl_ram_n_822, ZN => gl_ram_n_840);
  gl_ram_g9181 : ND2D0BWP7T port map(A1 => gl_ram_n_829, A2 => gl_ram_n_827, ZN => gl_ram_n_839);
  gl_ram_g9182 : ND2D0BWP7T port map(A1 => gl_ram_n_827, A2 => gl_ram_n_821, ZN => gl_ram_n_838);
  gl_ram_g9183 : ND2D0BWP7T port map(A1 => gl_ram_n_825, A2 => gl_ram_n_827, ZN => gl_ram_n_837);
  gl_ram_g9184 : ND2D0BWP7T port map(A1 => gl_ram_n_820, A2 => gl_ram_n_829, ZN => gl_ram_n_836);
  gl_ram_g9185 : OR2D1BWP7T port map(A1 => gl_ram_n_832, A2 => gl_ram_ram_position(1), Z => gl_ram_n_835);
  gl_ram_g9186 : CKND2D1BWP7T port map(A1 => gl_ram_n_830, A2 => gl_ram_ram_position(1), ZN => gl_ram_n_834);
  gl_ram_g9187 : CKND2D1BWP7T port map(A1 => gl_ram_n_831, A2 => gl_ram_ram_position(1), ZN => gl_ram_n_833);
  gl_ram_g9188 : ND2D0BWP7T port map(A1 => gl_ram_ram_position(2), A2 => gl_ram_ram_position(0), ZN => gl_ram_n_832);
  gl_ram_g9189 : NR2XD0BWP7T port map(A1 => FE_PHN505_sig_logic_x_0, A2 => sig_logic_x(1), ZN => gl_ram_n_1311);
  gl_ram_g9190 : NR2D0BWP7T port map(A1 => gl_ram_ram_position(0), A2 => gl_ram_ram_position(2), ZN => gl_ram_n_831);
  gl_ram_g9191 : INR2D0BWP7T port map(A1 => gl_ram_ram_position(2), B1 => gl_ram_ram_position(0), ZN => gl_ram_n_830);
  gl_ram_g9192 : INR2D0BWP7T port map(A1 => gl_ram_ram_position(4), B1 => gl_ram_ram_position(3), ZN => gl_ram_n_829);
  gl_ram_g9193 : ND2D0BWP7T port map(A1 => gl_ram_ram_position(3), A2 => gl_ram_ram_position(4), ZN => gl_ram_n_828);
  gl_ram_g9194 : INR2D0BWP7T port map(A1 => gl_ram_ram_position(6), B1 => gl_ram_ram_position(5), ZN => gl_ram_n_827);
  gl_ram_g9195 : INVD1BWP7T port map(I => gl_ram_n_823, ZN => gl_ram_n_824);
  gl_ram_g9196 : CKND2D0BWP7T port map(A1 => FE_PHN517_sig_logic_y_1, A2 => FE_PHN530_sig_logic_y_2, ZN => gl_ram_n_819);
  gl_ram_g9197 : INR2D0BWP7T port map(A1 => gl_ram_ram_position(0), B1 => gl_ram_ram_position(2), ZN => gl_ram_n_826);
  gl_ram_g9198 : INR2D0BWP7T port map(A1 => gl_ram_ram_position(3), B1 => gl_ram_ram_position(4), ZN => gl_ram_n_825);
  gl_ram_g9199 : ND2D1BWP7T port map(A1 => gl_sig_y(0), A2 => gl_sig_x(1), ZN => gl_ram_n_823);
  gl_ram_g9200 : NR2D0BWP7T port map(A1 => gl_ram_ram_position(5), A2 => gl_ram_ram_position(6), ZN => gl_ram_n_822);
  gl_ram_g9201 : NR2D0BWP7T port map(A1 => gl_ram_ram_position(4), A2 => gl_ram_ram_position(3), ZN => gl_ram_n_821);
  gl_ram_g9202 : INR2D0BWP7T port map(A1 => gl_ram_ram_position(5), B1 => gl_ram_ram_position(6), ZN => gl_ram_n_820);
  gl_ram_g9203 : CKND1BWP7T port map(I => FE_PHN516_sig_logic_y_3, ZN => gl_ram_n_1310);
  gl_ram_g2 : CKAN2D1BWP7T port map(A1 => gl_ram_n_1073, A2 => gl_ram_n_874, Z => gl_ram_n_818);
  gl_ram_ram_position_reg_0 : LHQD1BWP7T port map(D => gl_ram_x_grid(0), E => gl_ram_n_1111, Q => gl_ram_ram_position(0));
  gl_ram_ram_position_reg_1 : LHQD1BWP7T port map(D => gl_ram_n_407, E => gl_ram_n_1111, Q => gl_ram_ram_position(1));
  gl_ram_ram_position_reg_2 : LHQD1BWP7T port map(D => gl_ram_n_663, E => gl_ram_n_1111, Q => gl_ram_ram_position(2));
  gl_ram_ram_position_reg_3 : LHQD1BWP7T port map(D => gl_ram_n_730, E => gl_ram_n_1111, Q => gl_ram_ram_position(3));
  gl_ram_ram_position_reg_4 : LHQD1BWP7T port map(D => gl_ram_n_814, E => gl_ram_n_1111, Q => gl_ram_ram_position(4));
  gl_ram_ram_position_reg_5 : LHQD1BWP7T port map(D => gl_ram_n_815, E => gl_ram_n_1111, Q => gl_ram_ram_position(5));
  gl_ram_ram_position_reg_6 : LHQD1BWP7T port map(D => gl_ram_n_817, E => gl_ram_n_1111, Q => gl_ram_ram_position(6));
  gl_ram_ram_reg_0_0 : LNQD1BWP7T port map(D => gl_ram_n_1436, EN => gl_ram_n_812, Q => gl_ram_ram_0(0));
  gl_ram_ram_reg_0_1 : LNQD1BWP7T port map(D => gl_ram_n_1447, EN => gl_ram_n_812, Q => gl_ram_ram_0(1));
  gl_ram_ram_reg_0_2 : LNQD1BWP7T port map(D => gl_ram_n_1449, EN => gl_ram_n_812, Q => gl_ram_ram_0(2));
  gl_ram_ram_reg_1_0 : LNQD1BWP7T port map(D => gl_ram_n_736, EN => gl_ram_n_811, Q => gl_ram_ram_1(0));
  gl_ram_ram_reg_1_1 : LNQD1BWP7T port map(D => gl_ram_n_1447, EN => gl_ram_n_811, Q => gl_ram_ram_1(1));
  gl_ram_ram_reg_1_2 : LNQD1BWP7T port map(D => gl_ram_n_1449, EN => gl_ram_n_811, Q => gl_ram_ram_1(2));
  gl_ram_ram_reg_2_0 : LNQD1BWP7T port map(D => gl_ram_n_736, EN => gl_ram_n_810, Q => gl_ram_ram_2(0));
  gl_ram_ram_reg_2_1 : LNQD1BWP7T port map(D => gl_ram_n_1447, EN => gl_ram_n_810, Q => gl_ram_ram_2(1));
  gl_ram_ram_reg_2_2 : LNQD1BWP7T port map(D => gl_ram_n_1449, EN => gl_ram_n_810, Q => gl_ram_ram_2(2));
  gl_ram_ram_reg_3_0 : LNQD1BWP7T port map(D => gl_ram_n_736, EN => gl_ram_n_809, Q => gl_ram_ram_3(0));
  gl_ram_ram_reg_3_1 : LNQD1BWP7T port map(D => gl_ram_n_1446, EN => gl_ram_n_809, Q => gl_ram_ram_3(1));
  gl_ram_ram_reg_3_2 : LNQD2BWP7T port map(D => FE_OCPN1_gl_ram_n_1448, EN => gl_ram_n_809, Q => gl_ram_ram_3(2));
  gl_ram_ram_reg_4_0 : LNQD2BWP7T port map(D => gl_ram_n_736, EN => gl_ram_n_808, Q => gl_ram_ram_4(0));
  gl_ram_ram_reg_4_1 : LNQD1BWP7T port map(D => gl_ram_n_1446, EN => gl_ram_n_808, Q => gl_ram_ram_4(1));
  gl_ram_ram_reg_4_2 : LNQD2BWP7T port map(D => FE_OCPN1_gl_ram_n_1448, EN => gl_ram_n_808, Q => gl_ram_ram_4(2));
  gl_ram_ram_reg_5_0 : LNQD2BWP7T port map(D => gl_ram_n_736, EN => gl_ram_n_807, Q => gl_ram_ram_5(0));
  gl_ram_ram_reg_5_1 : LNQD1BWP7T port map(D => gl_ram_n_1446, EN => gl_ram_n_807, Q => gl_ram_ram_5(1));
  gl_ram_ram_reg_5_2 : LNQD1BWP7T port map(D => FE_OCPN1_gl_ram_n_1448, EN => gl_ram_n_807, Q => gl_ram_ram_5(2));
  gl_ram_ram_reg_6_0 : LNQD2BWP7T port map(D => gl_ram_n_736, EN => gl_ram_n_806, Q => gl_ram_ram_6(0));
  gl_ram_ram_reg_6_1 : LNQD1BWP7T port map(D => gl_ram_n_1446, EN => gl_ram_n_806, Q => gl_ram_ram_6(1));
  gl_ram_ram_reg_6_2 : LNQD1BWP7T port map(D => FE_OCPN1_gl_ram_n_1448, EN => gl_ram_n_806, Q => gl_ram_ram_6(2));
  gl_ram_ram_reg_7_0 : LNQD2BWP7T port map(D => gl_ram_n_736, EN => gl_ram_n_805, Q => gl_ram_ram_7(0));
  gl_ram_ram_reg_7_1 : LNQD1BWP7T port map(D => gl_ram_n_1447, EN => gl_ram_n_805, Q => gl_ram_ram_7(1));
  gl_ram_ram_reg_7_2 : LNQD1BWP7T port map(D => gl_ram_n_1449, EN => gl_ram_n_805, Q => gl_ram_ram_7(2));
  gl_ram_ram_reg_8_0 : LNQD1BWP7T port map(D => gl_ram_n_736, EN => gl_ram_n_804, Q => gl_ram_ram_8(0));
  gl_ram_ram_reg_8_1 : LNQD1BWP7T port map(D => gl_ram_n_1446, EN => gl_ram_n_804, Q => gl_ram_ram_8(1));
  gl_ram_ram_reg_8_2 : LNQD2BWP7T port map(D => FE_OCPN2_gl_ram_n_1448, EN => gl_ram_n_804, Q => gl_ram_ram_8(2));
  gl_ram_ram_reg_9_1 : LNQD1BWP7T port map(D => gl_ram_n_1446, EN => gl_ram_n_803, Q => gl_ram_ram_9(1));
  gl_ram_ram_reg_9_2 : LNQD2BWP7T port map(D => FE_OCPN2_gl_ram_n_1448, EN => gl_ram_n_803, Q => gl_ram_ram_9(2));
  gl_ram_ram_reg_10_0 : LNQD1BWP7T port map(D => gl_ram_n_736, EN => gl_ram_n_802, Q => gl_ram_ram_10(0));
  gl_ram_ram_reg_10_1 : LNQD1BWP7T port map(D => gl_ram_n_1447, EN => gl_ram_n_802, Q => gl_ram_ram_10(1));
  gl_ram_ram_reg_10_2 : LNQD1BWP7T port map(D => FE_OCPN2_gl_ram_n_1448, EN => gl_ram_n_802, Q => gl_ram_ram_10(2));
  gl_ram_ram_reg_11_0 : LNQD2BWP7T port map(D => gl_ram_n_736, EN => gl_ram_n_801, Q => gl_ram_ram_11(0));
  gl_ram_ram_reg_11_1 : LNQD1BWP7T port map(D => gl_ram_n_1446, EN => gl_ram_n_801, Q => gl_ram_ram_11(1));
  gl_ram_ram_reg_11_2 : LNQD2BWP7T port map(D => FE_OCPN2_gl_ram_n_1448, EN => gl_ram_n_801, Q => gl_ram_ram_11(2));
  gl_ram_ram_reg_12_1 : LNQD1BWP7T port map(D => gl_ram_n_1446, EN => gl_ram_n_800, Q => gl_ram_ram_12(1));
  gl_ram_ram_reg_12_2 : LNQD1BWP7T port map(D => FE_OCPN2_gl_ram_n_1448, EN => gl_ram_n_800, Q => gl_ram_ram_12(2));
  gl_ram_ram_reg_13_0 : LNQD1BWP7T port map(D => gl_ram_n_736, EN => gl_ram_n_799, Q => gl_ram_ram_13(0));
  gl_ram_ram_reg_13_1 : LNQD1BWP7T port map(D => gl_ram_n_1446, EN => gl_ram_n_799, Q => gl_ram_ram_13(1));
  gl_ram_ram_reg_13_2 : LNQD2BWP7T port map(D => FE_OCPN2_gl_ram_n_1448, EN => gl_ram_n_799, Q => gl_ram_ram_13(2));
  gl_ram_ram_reg_14_0 : LNQD1BWP7T port map(D => gl_ram_n_736, EN => gl_ram_n_798, Q => gl_ram_ram_14(0));
  gl_ram_ram_reg_14_1 : LNQD1BWP7T port map(D => gl_ram_n_1446, EN => gl_ram_n_798, Q => gl_ram_ram_14(1));
  gl_ram_ram_reg_14_2 : LNQD1BWP7T port map(D => FE_OCPN2_gl_ram_n_1448, EN => gl_ram_n_798, Q => gl_ram_ram_14(2));
  gl_ram_ram_reg_15_0 : LNQD1BWP7T port map(D => gl_ram_n_736, EN => gl_ram_n_797, Q => gl_ram_ram_15(0));
  gl_ram_ram_reg_15_1 : LNQD1BWP7T port map(D => gl_ram_n_1446, EN => gl_ram_n_797, Q => gl_ram_ram_15(1));
  gl_ram_ram_reg_15_2 : LNQD2BWP7T port map(D => FE_OCPN2_gl_ram_n_1448, EN => gl_ram_n_797, Q => gl_ram_ram_15(2));
  gl_ram_ram_reg_16_0 : LNQD1BWP7T port map(D => gl_ram_n_736, EN => gl_ram_n_796, Q => gl_ram_ram_16(0));
  gl_ram_ram_reg_16_1 : LNQD1BWP7T port map(D => gl_ram_n_1446, EN => gl_ram_n_796, Q => gl_ram_ram_16(1));
  gl_ram_ram_reg_16_2 : LNQD2BWP7T port map(D => FE_OCPN1_gl_ram_n_1448, EN => gl_ram_n_796, Q => gl_ram_ram_16(2));
  gl_ram_ram_reg_17_1 : LNQD1BWP7T port map(D => gl_ram_n_1446, EN => gl_ram_n_795, Q => gl_ram_ram_17(1));
  gl_ram_ram_reg_17_2 : LNQD1BWP7T port map(D => FE_OCPN1_gl_ram_n_1448, EN => gl_ram_n_795, Q => gl_ram_ram_17(2));
  gl_ram_ram_reg_18_0 : LNQD1BWP7T port map(D => gl_ram_n_736, EN => gl_ram_n_794, Q => gl_ram_ram_18(0));
  gl_ram_ram_reg_18_1 : LNQD1BWP7T port map(D => gl_ram_n_1446, EN => gl_ram_n_794, Q => gl_ram_ram_18(1));
  gl_ram_ram_reg_18_2 : LNQD1BWP7T port map(D => gl_ram_n_1449, EN => gl_ram_n_794, Q => gl_ram_ram_18(2));
  gl_ram_ram_reg_19_0 : LNQD1BWP7T port map(D => gl_ram_n_736, EN => gl_ram_n_793, Q => gl_ram_ram_19(0));
  gl_ram_ram_reg_19_1 : LNQD1BWP7T port map(D => gl_ram_n_1447, EN => gl_ram_n_793, Q => gl_ram_ram_19(1));
  gl_ram_ram_reg_19_2 : LNQD2BWP7T port map(D => gl_ram_n_1449, EN => gl_ram_n_793, Q => gl_ram_ram_19(2));
  gl_ram_ram_reg_20_0 : LNQD1BWP7T port map(D => gl_ram_n_736, EN => gl_ram_n_792, Q => gl_ram_ram_20(0));
  gl_ram_ram_reg_20_1 : LNQD1BWP7T port map(D => gl_ram_n_1447, EN => gl_ram_n_792, Q => gl_ram_ram_20(1));
  gl_ram_ram_reg_20_2 : LNQD1BWP7T port map(D => FE_OCPN2_gl_ram_n_1448, EN => gl_ram_n_792, Q => gl_ram_ram_20(2));
  gl_ram_ram_reg_21_0 : LNQD1BWP7T port map(D => gl_ram_n_736, EN => gl_ram_n_791, Q => gl_ram_ram_21(0));
  gl_ram_ram_reg_21_1 : LNQD1BWP7T port map(D => gl_ram_n_1446, EN => gl_ram_n_791, Q => gl_ram_ram_21(1));
  gl_ram_ram_reg_21_2 : LNQD1BWP7T port map(D => gl_ram_n_1449, EN => gl_ram_n_791, Q => gl_ram_ram_21(2));
  gl_ram_ram_reg_22_0 : LNQD1BWP7T port map(D => gl_ram_n_736, EN => gl_ram_n_790, Q => gl_ram_ram_22(0));
  gl_ram_ram_reg_22_1 : LNQD1BWP7T port map(D => gl_ram_n_1447, EN => gl_ram_n_790, Q => gl_ram_ram_22(1));
  gl_ram_ram_reg_22_2 : LNQD1BWP7T port map(D => FE_OCPN2_gl_ram_n_1448, EN => gl_ram_n_790, Q => gl_ram_ram_22(2));
  gl_ram_ram_reg_23_0 : LNQD1BWP7T port map(D => gl_ram_n_736, EN => gl_ram_n_789, Q => gl_ram_ram_23(0));
  gl_ram_ram_reg_23_1 : LNQD1BWP7T port map(D => gl_ram_n_1446, EN => gl_ram_n_789, Q => gl_ram_ram_23(1));
  gl_ram_ram_reg_23_2 : LNQD1BWP7T port map(D => gl_ram_n_1449, EN => gl_ram_n_789, Q => gl_ram_ram_23(2));
  gl_ram_ram_reg_24_0 : LNQD1BWP7T port map(D => gl_ram_n_1436, EN => gl_ram_n_788, Q => gl_ram_ram_24(0));
  gl_ram_ram_reg_24_1 : LNQD1BWP7T port map(D => gl_ram_n_1447, EN => gl_ram_n_788, Q => gl_ram_ram_24(1));
  gl_ram_ram_reg_24_2 : LNQD1BWP7T port map(D => gl_ram_n_1449, EN => gl_ram_n_788, Q => gl_ram_ram_24(2));
  gl_ram_ram_reg_25_1 : LNQD1BWP7T port map(D => gl_ram_n_1447, EN => gl_ram_n_787, Q => gl_ram_ram_25(1));
  gl_ram_ram_reg_25_2 : LNQD1BWP7T port map(D => gl_ram_n_1449, EN => gl_ram_n_787, Q => gl_ram_ram_25(2));
  gl_ram_ram_reg_26_1 : LNQD1BWP7T port map(D => gl_ram_n_1447, EN => gl_ram_n_786, Q => gl_ram_ram_26(1));
  gl_ram_ram_reg_26_2 : LNQD1BWP7T port map(D => gl_ram_n_1449, EN => gl_ram_n_786, Q => gl_ram_ram_26(2));
  gl_ram_ram_reg_27_0 : LNQD1BWP7T port map(D => gl_ram_n_1437, EN => gl_ram_n_785, Q => gl_ram_ram_27(0));
  gl_ram_ram_reg_27_1 : LNQD1BWP7T port map(D => gl_ram_n_1447, EN => gl_ram_n_785, Q => gl_ram_ram_27(1));
  gl_ram_ram_reg_27_2 : LNQD1BWP7T port map(D => gl_ram_n_1449, EN => gl_ram_n_785, Q => gl_ram_ram_27(2));
  gl_ram_ram_reg_29_0 : LNQD1BWP7T port map(D => gl_ram_n_1437, EN => gl_ram_n_783, Q => gl_ram_ram_29(0));
  gl_ram_ram_reg_29_1 : LNQD1BWP7T port map(D => gl_ram_n_1447, EN => gl_ram_n_783, Q => gl_ram_ram_29(1));
  gl_ram_ram_reg_29_2 : LNQD2BWP7T port map(D => gl_ram_n_1449, EN => gl_ram_n_783, Q => gl_ram_ram_29(2));
  gl_ram_ram_reg_31_0 : LNQD1BWP7T port map(D => gl_ram_n_1436, EN => gl_ram_n_781, Q => gl_ram_ram_31(0));
  gl_ram_ram_reg_32_0 : LNQD2BWP7T port map(D => gl_ram_n_1437, EN => gl_ram_n_780, Q => gl_ram_ram_32(0));
  gl_ram_ram_reg_32_1 : LNQD1BWP7T port map(D => gl_ram_n_1446, EN => gl_ram_n_780, Q => gl_ram_ram_32(1));
  gl_ram_ram_reg_32_2 : LNQD1BWP7T port map(D => gl_ram_n_1449, EN => gl_ram_n_780, Q => gl_ram_ram_32(2));
  gl_ram_ram_reg_33_1 : LNQD1BWP7T port map(D => gl_ram_n_1447, EN => gl_ram_n_779, Q => gl_ram_ram_33(1));
  gl_ram_ram_reg_33_2 : LNQD2BWP7T port map(D => FE_OCPN3_gl_ram_n_1448, EN => gl_ram_n_779, Q => gl_ram_ram_33(2));
  gl_ram_ram_reg_34_0 : LNQD1BWP7T port map(D => gl_ram_n_1437, EN => gl_ram_n_778, Q => gl_ram_ram_34(0));
  gl_ram_ram_reg_34_1 : LNQD1BWP7T port map(D => gl_ram_n_1446, EN => gl_ram_n_778, Q => gl_ram_ram_34(1));
  gl_ram_ram_reg_34_2 : LNQD2BWP7T port map(D => gl_ram_n_1449, EN => gl_ram_n_778, Q => gl_ram_ram_34(2));
  gl_ram_ram_reg_35_0 : LNQD2BWP7T port map(D => gl_ram_n_1437, EN => gl_ram_n_777, Q => gl_ram_ram_35(0));
  gl_ram_ram_reg_35_1 : LNQD1BWP7T port map(D => gl_ram_n_1447, EN => gl_ram_n_777, Q => gl_ram_ram_35(1));
  gl_ram_ram_reg_35_2 : LNQD2BWP7T port map(D => gl_ram_n_1449, EN => gl_ram_n_777, Q => gl_ram_ram_35(2));
  gl_ram_ram_reg_36_0 : LNQD1BWP7T port map(D => gl_ram_n_1437, EN => gl_ram_n_776, Q => gl_ram_ram_36(0));
  gl_ram_ram_reg_36_1 : LNQD1BWP7T port map(D => gl_ram_n_1447, EN => gl_ram_n_776, Q => gl_ram_ram_36(1));
  gl_ram_ram_reg_36_2 : LNQD2BWP7T port map(D => FE_OCPN3_gl_ram_n_1448, EN => gl_ram_n_776, Q => gl_ram_ram_36(2));
  gl_ram_ram_reg_37_0 : LNQD1BWP7T port map(D => gl_ram_n_1437, EN => gl_ram_n_775, Q => gl_ram_ram_37(0));
  gl_ram_ram_reg_37_1 : LNQD1BWP7T port map(D => gl_ram_n_1446, EN => gl_ram_n_775, Q => gl_ram_ram_37(1));
  gl_ram_ram_reg_37_2 : LNQD1BWP7T port map(D => gl_ram_n_1449, EN => gl_ram_n_775, Q => gl_ram_ram_37(2));
  gl_ram_ram_reg_38_0 : LNQD1BWP7T port map(D => gl_ram_n_1437, EN => gl_ram_n_774, Q => gl_ram_ram_38(0));
  gl_ram_ram_reg_38_1 : LNQD1BWP7T port map(D => gl_ram_n_1447, EN => gl_ram_n_774, Q => gl_ram_ram_38(1));
  gl_ram_ram_reg_38_2 : LNQD1BWP7T port map(D => gl_ram_n_1449, EN => gl_ram_n_774, Q => gl_ram_ram_38(2));
  gl_ram_ram_reg_39_0 : LNQD1BWP7T port map(D => gl_ram_n_1437, EN => gl_ram_n_773, Q => gl_ram_ram_39(0));
  gl_ram_ram_reg_39_1 : LNQD1BWP7T port map(D => gl_ram_n_1447, EN => gl_ram_n_773, Q => gl_ram_ram_39(1));
  gl_ram_ram_reg_39_2 : LNQD2BWP7T port map(D => FE_OCPN3_gl_ram_n_1448, EN => gl_ram_n_773, Q => gl_ram_ram_39(2));
  gl_ram_ram_reg_40_0 : LNQD2BWP7T port map(D => gl_ram_n_1437, EN => gl_ram_n_772, Q => gl_ram_ram_40(0));
  gl_ram_ram_reg_40_1 : LNQD1BWP7T port map(D => gl_ram_n_1446, EN => gl_ram_n_772, Q => gl_ram_ram_40(1));
  gl_ram_ram_reg_40_2 : LNQD1BWP7T port map(D => gl_ram_n_1449, EN => gl_ram_n_772, Q => gl_ram_ram_40(2));
  gl_ram_ram_reg_42_0 : LNQD1BWP7T port map(D => gl_ram_n_1437, EN => gl_ram_n_770, Q => gl_ram_ram_42(0));
  gl_ram_ram_reg_42_1 : LNQD1BWP7T port map(D => gl_ram_n_1446, EN => gl_ram_n_770, Q => gl_ram_ram_42(1));
  gl_ram_ram_reg_42_2 : LNQD1BWP7T port map(D => gl_ram_n_1449, EN => gl_ram_n_770, Q => gl_ram_ram_42(2));
  gl_ram_ram_reg_43_0 : LNQD2BWP7T port map(D => gl_ram_n_1436, EN => gl_ram_n_769, Q => gl_ram_ram_43(0));
  gl_ram_ram_reg_43_1 : LNQD1BWP7T port map(D => gl_ram_n_1446, EN => gl_ram_n_769, Q => gl_ram_ram_43(1));
  gl_ram_ram_reg_43_2 : LNQD2BWP7T port map(D => FE_OCPN3_gl_ram_n_1448, EN => gl_ram_n_769, Q => gl_ram_ram_43(2));
  gl_ram_ram_reg_44_0 : LNQD1BWP7T port map(D => gl_ram_n_1436, EN => gl_ram_n_768, Q => gl_ram_ram_44(0));
  gl_ram_ram_reg_44_1 : LNQD1BWP7T port map(D => gl_ram_n_1447, EN => gl_ram_n_768, Q => gl_ram_ram_44(1));
  gl_ram_ram_reg_44_2 : LNQD1BWP7T port map(D => gl_ram_n_1449, EN => gl_ram_n_768, Q => gl_ram_ram_44(2));
  gl_ram_ram_reg_45_0 : LNQD1BWP7T port map(D => gl_ram_n_1437, EN => gl_ram_n_767, Q => gl_ram_ram_45(0));
  gl_ram_ram_reg_45_1 : LNQD1BWP7T port map(D => gl_ram_n_1446, EN => gl_ram_n_767, Q => gl_ram_ram_45(1));
  gl_ram_ram_reg_45_2 : LNQD1BWP7T port map(D => gl_ram_n_1449, EN => gl_ram_n_767, Q => gl_ram_ram_45(2));
  gl_ram_ram_reg_46_0 : LNQD2BWP7T port map(D => gl_ram_n_1437, EN => gl_ram_n_766, Q => gl_ram_ram_46(0));
  gl_ram_ram_reg_46_1 : LNQD1BWP7T port map(D => gl_ram_n_1447, EN => gl_ram_n_766, Q => gl_ram_ram_46(1));
  gl_ram_ram_reg_46_2 : LNQD1BWP7T port map(D => gl_ram_n_1449, EN => gl_ram_n_766, Q => gl_ram_ram_46(2));
  gl_ram_ram_reg_47_0 : LNQD1BWP7T port map(D => gl_ram_n_1436, EN => gl_ram_n_765, Q => gl_ram_ram_47(0));
  gl_ram_ram_reg_47_1 : LNQD1BWP7T port map(D => gl_ram_n_1447, EN => gl_ram_n_765, Q => gl_ram_ram_47(1));
  gl_ram_ram_reg_47_2 : LNQD1BWP7T port map(D => gl_ram_n_1449, EN => gl_ram_n_765, Q => gl_ram_ram_47(2));
  gl_ram_ram_reg_48_0 : LNQD2BWP7T port map(D => gl_ram_n_1436, EN => gl_ram_n_764, Q => gl_ram_ram_48(0));
  gl_ram_ram_reg_48_1 : LNQD1BWP7T port map(D => gl_ram_n_1447, EN => gl_ram_n_764, Q => gl_ram_ram_48(1));
  gl_ram_ram_reg_48_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => gl_ram_n_764, Q => gl_ram_ram_48(2));
  gl_ram_ram_reg_49_0 : LNQD2BWP7T port map(D => gl_ram_n_1436, EN => gl_ram_n_763, Q => gl_ram_ram_49(0));
  gl_ram_ram_reg_49_1 : LNQD1BWP7T port map(D => gl_ram_n_1447, EN => gl_ram_n_763, Q => gl_ram_ram_49(1));
  gl_ram_ram_reg_49_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => gl_ram_n_763, Q => gl_ram_ram_49(2));
  gl_ram_ram_reg_50_0 : LNQD2BWP7T port map(D => gl_ram_n_1436, EN => gl_ram_n_762, Q => gl_ram_ram_50(0));
  gl_ram_ram_reg_50_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => gl_ram_n_762, Q => gl_ram_ram_50(1));
  gl_ram_ram_reg_50_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => gl_ram_n_762, Q => gl_ram_ram_50(2));
  gl_ram_ram_reg_51_0 : LNQD2BWP7T port map(D => gl_ram_n_1436, EN => gl_ram_n_761, Q => gl_ram_ram_51(0));
  gl_ram_ram_reg_51_1 : LNQD2BWP7T port map(D => gl_ram_n_735, EN => gl_ram_n_761, Q => gl_ram_ram_51(1));
  gl_ram_ram_reg_51_2 : LNQD2BWP7T port map(D => gl_ram_n_739, EN => gl_ram_n_761, Q => gl_ram_ram_51(2));
  gl_ram_ram_reg_52_0 : LNQD2BWP7T port map(D => gl_ram_n_1436, EN => gl_ram_n_760, Q => gl_ram_ram_52(0));
  gl_ram_ram_reg_52_1 : LNQD2BWP7T port map(D => gl_ram_n_735, EN => gl_ram_n_760, Q => gl_ram_ram_52(1));
  gl_ram_ram_reg_52_2 : LNQD2BWP7T port map(D => gl_ram_n_739, EN => gl_ram_n_760, Q => gl_ram_ram_52(2));
  gl_ram_ram_reg_53_0 : LNQD2BWP7T port map(D => gl_ram_n_1436, EN => gl_ram_n_759, Q => gl_ram_ram_53(0));
  gl_ram_ram_reg_53_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => gl_ram_n_759, Q => gl_ram_ram_53(1));
  gl_ram_ram_reg_53_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => gl_ram_n_759, Q => gl_ram_ram_53(2));
  gl_ram_ram_reg_54_0 : LNQD2BWP7T port map(D => gl_ram_n_1437, EN => gl_ram_n_758, Q => gl_ram_ram_54(0));
  gl_ram_ram_reg_54_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => gl_ram_n_758, Q => gl_ram_ram_54(1));
  gl_ram_ram_reg_54_2 : LNQD2BWP7T port map(D => gl_ram_n_739, EN => gl_ram_n_758, Q => gl_ram_ram_54(2));
  gl_ram_ram_reg_55_0 : LNQD2BWP7T port map(D => gl_ram_n_1437, EN => gl_ram_n_757, Q => gl_ram_ram_55(0));
  gl_ram_ram_reg_55_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => gl_ram_n_757, Q => gl_ram_ram_55(1));
  gl_ram_ram_reg_55_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => gl_ram_n_757, Q => gl_ram_ram_55(2));
  gl_ram_ram_reg_56_0 : LNQD1BWP7T port map(D => gl_ram_n_1436, EN => gl_ram_n_756, Q => gl_ram_ram_56(0));
  gl_ram_ram_reg_56_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => gl_ram_n_756, Q => gl_ram_ram_56(1));
  gl_ram_ram_reg_56_2 : LNQD2BWP7T port map(D => gl_ram_n_739, EN => gl_ram_n_756, Q => gl_ram_ram_56(2));
  gl_ram_ram_reg_59_0 : LNQD1BWP7T port map(D => gl_ram_n_1436, EN => gl_ram_n_753, Q => gl_ram_ram_59(0));
  gl_ram_ram_reg_59_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => gl_ram_n_753, Q => gl_ram_ram_59(1));
  gl_ram_ram_reg_59_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => gl_ram_n_753, Q => gl_ram_ram_59(2));
  gl_ram_ram_reg_60_0 : LNQD1BWP7T port map(D => gl_ram_n_1437, EN => gl_ram_n_752, Q => gl_ram_ram_60(0));
  gl_ram_ram_reg_60_1 : LNQD2BWP7T port map(D => gl_ram_n_735, EN => gl_ram_n_752, Q => gl_ram_ram_60(1));
  gl_ram_ram_reg_60_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => gl_ram_n_752, Q => gl_ram_ram_60(2));
  gl_ram_ram_reg_61_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => gl_ram_n_751, Q => gl_ram_ram_61(1));
  gl_ram_ram_reg_61_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => gl_ram_n_751, Q => gl_ram_ram_61(2));
  gl_ram_ram_reg_62_0 : LNQD1BWP7T port map(D => gl_ram_n_1436, EN => gl_ram_n_750, Q => gl_ram_ram_62(0));
  gl_ram_ram_reg_62_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => gl_ram_n_750, Q => gl_ram_ram_62(1));
  gl_ram_ram_reg_62_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => gl_ram_n_750, Q => gl_ram_ram_62(2));
  gl_ram_ram_reg_63_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => gl_ram_n_749, Q => gl_ram_ram_63(1));
  gl_ram_ram_reg_63_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => gl_ram_n_749, Q => gl_ram_ram_63(2));
  gl_ram_ram_reg_64_0 : LHCNQD2BWP7T port map(CDN => FE_OFN32_logic_1_1_net, D => gl_ram_n_736, E => CTS_306, Q => gl_ram_ram_64(0));
  gl_ram_ram_reg_64_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => CTS_307, Q => gl_ram_ram_64(1));
  gl_ram_ram_reg_64_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => CTS_307, Q => gl_ram_ram_64(2));
  gl_ram_ram_reg_65_0 : LHCNQD2BWP7T port map(CDN => FE_OFN32_logic_1_1_net, D => gl_ram_n_736, E => CTS_299, Q => gl_ram_ram_65(0));
  gl_ram_ram_reg_65_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => CTS_300, Q => gl_ram_ram_65(1));
  gl_ram_ram_reg_65_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => CTS_300, Q => gl_ram_ram_65(2));
  gl_ram_ram_reg_66_0 : LHCNQD2BWP7T port map(CDN => FE_OFN32_logic_1_1_net, D => gl_ram_n_736, E => CTS_302, Q => gl_ram_ram_66(0));
  gl_ram_ram_reg_66_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => CTS_303, Q => gl_ram_ram_66(1));
  gl_ram_ram_reg_66_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => CTS_303, Q => gl_ram_ram_66(2));
  gl_ram_ram_reg_67_0 : LHCNQD2BWP7T port map(CDN => FE_OFN32_logic_1_1_net, D => gl_ram_n_736, E => CTS_309, Q => gl_ram_ram_67(0));
  gl_ram_ram_reg_67_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => CTS_310, Q => gl_ram_ram_67(1));
  gl_ram_ram_reg_67_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => CTS_310, Q => gl_ram_ram_67(2));
  gl_ram_ram_reg_68_0 : LHCNQD2BWP7T port map(CDN => FE_OFN32_logic_1_1_net, D => gl_ram_n_736, E => CTS_358, Q => gl_ram_ram_68(0));
  gl_ram_ram_reg_68_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => CTS_359, Q => gl_ram_ram_68(1));
  gl_ram_ram_reg_68_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => CTS_359, Q => gl_ram_ram_68(2));
  gl_ram_ram_reg_69_0 : LHCNQD2BWP7T port map(CDN => FE_OFN32_logic_1_1_net, D => gl_ram_n_736, E => CTS_355, Q => gl_ram_ram_69(0));
  gl_ram_ram_reg_69_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => CTS_356, Q => gl_ram_ram_69(1));
  gl_ram_ram_reg_69_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => CTS_356, Q => gl_ram_ram_69(2));
  gl_ram_ram_reg_70_0 : LHCNQD1BWP7T port map(CDN => FE_OFN32_logic_1_1_net, D => gl_ram_n_736, E => CTS_285, Q => gl_ram_ram_70(0));
  gl_ram_ram_reg_70_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => CTS_286, Q => gl_ram_ram_70(1));
  gl_ram_ram_reg_70_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => CTS_286, Q => gl_ram_ram_70(2));
  gl_ram_ram_reg_71_0 : LHCNQD2BWP7T port map(CDN => FE_OFN32_logic_1_1_net, D => gl_ram_n_736, E => CTS_361, Q => gl_ram_ram_71(0));
  gl_ram_ram_reg_71_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => CTS_362, Q => gl_ram_ram_71(1));
  gl_ram_ram_reg_71_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => CTS_362, Q => gl_ram_ram_71(2));
  gl_ram_ram_reg_72_0 : LHCNQD2BWP7T port map(CDN => FE_OFN32_logic_1_1_net, D => gl_ram_n_736, E => CTS_332, Q => gl_ram_ram_72(0));
  gl_ram_ram_reg_72_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => CTS_333, Q => gl_ram_ram_72(1));
  gl_ram_ram_reg_72_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => CTS_333, Q => gl_ram_ram_72(2));
  gl_ram_ram_reg_73_0 : LHCNQD2BWP7T port map(CDN => FE_OFN32_logic_1_1_net, D => gl_ram_n_736, E => CTS_334, Q => gl_ram_ram_73(0));
  gl_ram_ram_reg_73_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => CTS_335, Q => gl_ram_ram_73(1));
  gl_ram_ram_reg_73_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => CTS_335, Q => gl_ram_ram_73(2));
  gl_ram_ram_reg_74_0 : LHCNQD2BWP7T port map(CDN => FE_OFN32_logic_1_1_net, D => gl_ram_n_736, E => CTS_297, Q => gl_ram_ram_74(0));
  gl_ram_ram_reg_74_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => CTS_298, Q => gl_ram_ram_74(1));
  gl_ram_ram_reg_74_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => CTS_298, Q => gl_ram_ram_74(2));
  gl_ram_ram_reg_75_0 : LHCNQD2BWP7T port map(CDN => FE_OFN32_logic_1_1_net, D => gl_ram_n_736, E => CTS_293, Q => gl_ram_ram_75(0));
  gl_ram_ram_reg_75_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => CTS_294, Q => gl_ram_ram_75(1));
  gl_ram_ram_reg_75_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => CTS_294, Q => gl_ram_ram_75(2));
  gl_ram_ram_reg_76_0 : LHCNQD2BWP7T port map(CDN => FE_OFN32_logic_1_1_net, D => gl_ram_n_736, E => CTS_340, Q => gl_ram_ram_76(0));
  gl_ram_ram_reg_76_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => CTS_341, Q => gl_ram_ram_76(1));
  gl_ram_ram_reg_76_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => CTS_341, Q => gl_ram_ram_76(2));
  gl_ram_ram_reg_77_0 : LNQD1BWP7T port map(D => gl_ram_n_1436, EN => gl_ram_n_748, Q => gl_ram_ram_77(0));
  gl_ram_ram_reg_77_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => gl_ram_n_748, Q => gl_ram_ram_77(1));
  gl_ram_ram_reg_77_2 : LNQD1BWP7T port map(D => FE_OCPN1_gl_ram_n_1448, EN => gl_ram_n_748, Q => gl_ram_ram_77(2));
  gl_ram_ram_reg_78_0 : LHCNQD2BWP7T port map(CDN => FE_OFN32_logic_1_1_net, D => gl_ram_n_736, E => CTS_312, Q => gl_ram_ram_78(0));
  gl_ram_ram_reg_78_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => CTS_313, Q => gl_ram_ram_78(1));
  gl_ram_ram_reg_78_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => CTS_313, Q => gl_ram_ram_78(2));
  gl_ram_ram_reg_79_0 : LHCNQD2BWP7T port map(CDN => FE_OFN32_logic_1_1_net, D => gl_ram_n_736, E => CTS_336, Q => gl_ram_ram_79(0));
  gl_ram_ram_reg_79_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => CTS_337, Q => gl_ram_ram_79(1));
  gl_ram_ram_reg_79_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => CTS_337, Q => gl_ram_ram_79(2));
  gl_ram_ram_reg_80_0 : LHCNQD2BWP7T port map(CDN => FE_OFN32_logic_1_1_net, D => gl_ram_n_736, E => CTS_290, Q => gl_ram_ram_80(0));
  gl_ram_ram_reg_80_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => CTS_291, Q => gl_ram_ram_80(1));
  gl_ram_ram_reg_80_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => CTS_291, Q => gl_ram_ram_80(2));
  gl_ram_ram_reg_81_0 : LHCNQD2BWP7T port map(CDN => FE_OFN32_logic_1_1_net, D => gl_ram_n_736, E => CTS_315, Q => gl_ram_ram_81(0));
  gl_ram_ram_reg_81_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => CTS_316, Q => gl_ram_ram_81(1));
  gl_ram_ram_reg_81_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => CTS_316, Q => gl_ram_ram_81(2));
  gl_ram_ram_reg_82_0 : LHCNQD2BWP7T port map(CDN => FE_OFN32_logic_1_1_net, D => gl_ram_n_736, E => CTS_330, Q => gl_ram_ram_82(0));
  gl_ram_ram_reg_82_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => CTS_331, Q => gl_ram_ram_82(1));
  gl_ram_ram_reg_82_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => CTS_331, Q => gl_ram_ram_82(2));
  gl_ram_ram_reg_83_0 : LHCNQD2BWP7T port map(CDN => FE_OFN32_logic_1_1_net, D => gl_ram_n_736, E => CTS_338, Q => gl_ram_ram_83(0));
  gl_ram_ram_reg_83_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => CTS_339, Q => gl_ram_ram_83(1));
  gl_ram_ram_reg_83_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => CTS_339, Q => gl_ram_ram_83(2));
  gl_ram_ram_reg_84_0 : LHCNQD2BWP7T port map(CDN => FE_OFN32_logic_1_1_net, D => gl_ram_n_736, E => CTS_346, Q => gl_ram_ram_84(0));
  gl_ram_ram_reg_84_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => CTS_347, Q => gl_ram_ram_84(1));
  gl_ram_ram_reg_84_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => CTS_347, Q => gl_ram_ram_84(2));
  gl_ram_ram_reg_85_0 : LHCNQD2BWP7T port map(CDN => FE_OFN32_logic_1_1_net, D => gl_ram_n_736, E => CTS_324, Q => gl_ram_ram_85(0));
  gl_ram_ram_reg_85_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => CTS_325, Q => gl_ram_ram_85(1));
  gl_ram_ram_reg_85_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => CTS_325, Q => gl_ram_ram_85(2));
  gl_ram_ram_reg_86_0 : LHCNQD2BWP7T port map(CDN => FE_OFN32_logic_1_1_net, D => gl_ram_n_736, E => CTS_328, Q => gl_ram_ram_86(0));
  gl_ram_ram_reg_86_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => CTS_329, Q => gl_ram_ram_86(1));
  gl_ram_ram_reg_86_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => CTS_329, Q => gl_ram_ram_86(2));
  gl_ram_ram_reg_87_0 : LHCNQD2BWP7T port map(CDN => FE_OFN32_logic_1_1_net, D => gl_ram_n_736, E => CTS_319, Q => gl_ram_ram_87(0));
  gl_ram_ram_reg_87_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => CTS_320, Q => gl_ram_ram_87(1));
  gl_ram_ram_reg_87_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => CTS_320, Q => gl_ram_ram_87(2));
  gl_ram_ram_reg_88_0 : LNQD1BWP7T port map(D => gl_ram_n_1437, EN => gl_ram_n_747, Q => gl_ram_ram_88(0));
  gl_ram_ram_reg_88_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => gl_ram_n_747, Q => gl_ram_ram_88(1));
  gl_ram_ram_reg_88_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => gl_ram_n_747, Q => gl_ram_ram_88(2));
  gl_ram_ram_reg_89_0 : LNQD1BWP7T port map(D => gl_ram_n_1437, EN => gl_ram_n_746, Q => gl_ram_ram_89(0));
  gl_ram_ram_reg_89_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => gl_ram_n_746, Q => gl_ram_ram_89(1));
  gl_ram_ram_reg_89_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => gl_ram_n_746, Q => gl_ram_ram_89(2));
  gl_ram_ram_reg_90_0 : LNQD1BWP7T port map(D => gl_ram_n_1436, EN => gl_ram_n_745, Q => gl_ram_ram_90(0));
  gl_ram_ram_reg_90_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => gl_ram_n_745, Q => gl_ram_ram_90(1));
  gl_ram_ram_reg_90_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => gl_ram_n_745, Q => gl_ram_ram_90(2));
  gl_ram_ram_reg_91_0 : LNQD1BWP7T port map(D => gl_ram_n_1437, EN => gl_ram_n_744, Q => gl_ram_ram_91(0));
  gl_ram_ram_reg_91_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => gl_ram_n_744, Q => gl_ram_ram_91(1));
  gl_ram_ram_reg_91_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => gl_ram_n_744, Q => gl_ram_ram_91(2));
  gl_ram_ram_reg_92_0 : LNQD1BWP7T port map(D => gl_ram_n_1436, EN => gl_ram_n_743, Q => gl_ram_ram_92(0));
  gl_ram_ram_reg_92_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => gl_ram_n_743, Q => gl_ram_ram_92(1));
  gl_ram_ram_reg_92_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => gl_ram_n_743, Q => gl_ram_ram_92(2));
  gl_ram_ram_reg_93_0 : LNQD1BWP7T port map(D => gl_ram_n_1436, EN => gl_ram_n_742, Q => gl_ram_ram_93(0));
  gl_ram_ram_reg_93_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => gl_ram_n_742, Q => gl_ram_ram_93(1));
  gl_ram_ram_reg_93_2 : LNQD1BWP7T port map(D => FE_OCPN2_gl_ram_n_1448, EN => gl_ram_n_742, Q => gl_ram_ram_93(2));
  gl_ram_ram_reg_94_0 : LNQD1BWP7T port map(D => gl_ram_n_1436, EN => gl_ram_n_741, Q => gl_ram_ram_94(0));
  gl_ram_ram_reg_94_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => gl_ram_n_741, Q => gl_ram_ram_94(1));
  gl_ram_ram_reg_94_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => gl_ram_n_741, Q => gl_ram_ram_94(2));
  gl_ram_ram_reg_95_0 : LNQD1BWP7T port map(D => gl_ram_n_1436, EN => gl_ram_n_740, Q => gl_ram_ram_95(0));
  gl_ram_ram_reg_95_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => gl_ram_n_740, Q => gl_ram_ram_95(1));
  gl_ram_ram_reg_95_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => gl_ram_n_740, Q => gl_ram_ram_95(2));
  gl_ram_ram_reg_96_0 : LHCNQD2BWP7T port map(CDN => FE_OFN32_logic_1_1_net, D => gl_ram_n_736, E => CTS_352, Q => gl_ram_ram_96(0));
  gl_ram_ram_reg_96_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => CTS_353, Q => gl_ram_ram_96(1));
  gl_ram_ram_reg_96_2 : LNQD2BWP7T port map(D => gl_ram_n_739, EN => CTS_353, Q => gl_ram_ram_96(2));
  gl_ram_ram_reg_97_0 : LHCNQD2BWP7T port map(CDN => FE_OFN32_logic_1_1_net, D => gl_ram_n_736, E => CTS_326, Q => gl_ram_ram_97(0));
  gl_ram_ram_reg_97_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => CTS_327, Q => gl_ram_ram_97(1));
  gl_ram_ram_reg_97_2 : LNQD2BWP7T port map(D => gl_ram_n_739, EN => CTS_327, Q => gl_ram_ram_97(2));
  gl_ram_ram_reg_98_0 : LHCNQD2BWP7T port map(CDN => FE_OFN32_logic_1_1_net, D => gl_ram_n_736, E => CTS_342, Q => gl_ram_ram_98(0));
  gl_ram_ram_reg_98_1 : LNQD2BWP7T port map(D => gl_ram_n_735, EN => CTS_343, Q => gl_ram_ram_98(1));
  gl_ram_ram_reg_98_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => CTS_343, Q => gl_ram_ram_98(2));
  gl_ram_ram_reg_99_0 : LHCNQD2BWP7T port map(CDN => FE_OFN32_logic_1_1_net, D => gl_ram_n_736, E => CTS_349, Q => gl_ram_ram_99(0));
  gl_ram_ram_reg_99_1 : LNQD1BWP7T port map(D => gl_ram_n_735, EN => CTS_350, Q => gl_ram_ram_99(1));
  gl_ram_ram_reg_99_2 : LNQD1BWP7T port map(D => gl_ram_n_739, EN => CTS_350, Q => gl_ram_ram_99(2));
  gl_ram_x_grid_reg_0 : LHQD1BWP7T port map(D => gl_ram_n_18, E => gl_ram_n_1111, Q => gl_ram_x_grid(0));
  gl_ram_x_grid_reg_1 : LHQD1BWP7T port map(D => gl_ram_n_34, E => gl_ram_n_1111, Q => gl_ram_x_grid(1));
  gl_ram_x_grid_reg_2 : LHQD1BWP7T port map(D => gl_ram_n_85, E => gl_ram_n_1111, Q => gl_ram_x_grid(2));
  gl_ram_x_grid_reg_3 : LHQD1BWP7T port map(D => gl_ram_n_572, E => gl_ram_n_1111, Q => gl_ram_x_grid(3));
  gl_ram_x_grid_reg_4 : LHQD1BWP7T port map(D => gl_ram_n_1320, E => gl_ram_n_1111, Q => gl_ram_x_grid(4));
  gl_ram_y_grid_reg_0 : LHQD1BWP7T port map(D => gl_ram_n_19, E => gl_ram_n_1111, Q => gl_ram_y_grid(0));
  gl_ram_y_grid_reg_1 : LHQD1BWP7T port map(D => gl_ram_n_35, E => gl_ram_n_1111, Q => gl_ram_y_grid(1));
  gl_ram_y_grid_reg_2 : LHQD1BWP7T port map(D => gl_ram_n_661, E => gl_ram_n_1111, Q => gl_ram_y_grid(2));
  gl_ram_y_grid_reg_3 : LHQD1BWP7T port map(D => gl_ram_n_698, E => gl_ram_n_1111, Q => gl_ram_y_grid(3));
  gl_ram_y_grid_reg_4 : LHQD1BWP7T port map(D => gl_ram_n_695, E => gl_ram_n_1111, Q => gl_ram_y_grid(4));
  gl_ram_g55626 : MOAI22D0BWP7T port map(A1 => gl_ram_n_816, A2 => gl_ram_n_679, B1 => gl_ram_n_816, B2 => gl_ram_n_679, ZN => gl_ram_n_817);
  gl_ram_g55628 : FA1D0BWP7T port map(A => gl_ram_n_410, B => gl_ram_n_652, CI => gl_ram_n_813, CO => gl_ram_n_816, S => gl_ram_n_815);
  gl_ram_g55630 : FA1D0BWP7T port map(A => gl_ram_n_653, B => gl_ram_n_404, CI => gl_ram_n_729, CO => gl_ram_n_813, S => gl_ram_n_814);
  gl_ram_g55932 : ND2D8BWP7T port map(A1 => gl_ram_n_733, A2 => gl_ram_n_728, ZN => gl_ram_n_739);
  gl_ram_g55935 : ND2D8BWP7T port map(A1 => gl_ram_n_732, A2 => gl_ram_n_727, ZN => gl_ram_n_736);
  gl_ram_g55936 : ND2D8BWP7T port map(A1 => gl_ram_n_731, A2 => gl_ram_n_726, ZN => gl_ram_n_735);
  gl_ram_g55938 : FA1D0BWP7T port map(A => gl_ram_n_405, B => gl_ram_y_grid(2), CI => gl_ram_n_662, CO => gl_ram_n_729, S => gl_ram_n_730);
  gl_ram_g55939 : ND2D6BWP7T port map(A1 => gl_ram_n_722, A2 => gl_ram_n_109, ZN => gl_ram_n_733);
  gl_ram_g55940 : ND2D8BWP7T port map(A1 => gl_ram_n_721, A2 => gl_ram_n_109, ZN => gl_ram_n_732);
  gl_ram_g55941 : ND2D6BWP7T port map(A1 => gl_ram_n_720, A2 => gl_ram_n_109, ZN => gl_ram_n_731);
  gl_ram_g55942 : NR2XD8BWP7T port map(A1 => gl_ram_n_725, A2 => gl_ram_n_701, ZN => gl_ram_n_728);
  gl_ram_g55943 : NR2XD8BWP7T port map(A1 => gl_ram_n_724, A2 => gl_ram_n_700, ZN => gl_ram_n_727);
  gl_ram_g55944 : NR2XD8BWP7T port map(A1 => gl_ram_n_723, A2 => gl_ram_n_699, ZN => gl_ram_n_726);
  gl_ram_g55945 : ND2D4BWP7T port map(A1 => gl_ram_n_719, A2 => gl_ram_n_1549, ZN => gl_ram_n_725);
  gl_ram_g55946 : ND2D6BWP7T port map(A1 => gl_ram_n_718, A2 => gl_ram_n_8, ZN => gl_ram_n_724);
  gl_ram_g55947 : ND2D4BWP7T port map(A1 => gl_ram_n_717, A2 => gl_ram_n_1550, ZN => gl_ram_n_723);
  gl_ram_g55948 : ND4D4BWP7T port map(A1 => gl_ram_n_712, A2 => gl_ram_n_709, A3 => gl_ram_n_710, A4 => gl_ram_n_716, ZN => gl_ram_n_722);
  gl_ram_g55949 : ND4D4BWP7T port map(A1 => gl_ram_n_711, A2 => gl_ram_n_705, A3 => gl_ram_n_707, A4 => gl_ram_n_706, ZN => gl_ram_n_721);
  gl_ram_g55951 : NR2XD2BWP7T port map(A1 => gl_ram_n_708, A2 => gl_ram_n_669, ZN => gl_ram_n_719);
  gl_ram_g55953 : NR2D4BWP7T port map(A1 => gl_ram_n_715, A2 => gl_ram_n_668, ZN => gl_ram_n_718);
  gl_ram_g55954 : NR2D4BWP7T port map(A1 => gl_ram_n_714, A2 => gl_ram_n_665, ZN => gl_ram_n_717);
  gl_ram_g55955 : NR2XD3BWP7T port map(A1 => gl_ram_n_687, A2 => gl_ram_n_682, ZN => gl_ram_n_716);
  gl_ram_g55956 : AOI21D2BWP7T port map(A1 => gl_ram_n_660, A2 => gl_ram_n_1451, B => gl_ram_n_409, ZN => gl_ram_n_715);
  gl_ram_g55958 : NR2XD2BWP7T port map(A1 => gl_ram_n_696, A2 => gl_ram_n_677, ZN => gl_ram_n_713);
  gl_ram_g55959 : NR2XD2BWP7T port map(A1 => gl_ram_n_694, A2 => gl_ram_n_675, ZN => gl_ram_n_712);
  gl_ram_g55960 : NR2XD3BWP7T port map(A1 => gl_ram_n_673, A2 => gl_ram_n_693, ZN => gl_ram_n_711);
  gl_ram_g55961 : NR2XD3BWP7T port map(A1 => gl_ram_n_692, A2 => gl_ram_n_676, ZN => gl_ram_n_710);
  gl_ram_g55962 : NR2XD3BWP7T port map(A1 => gl_ram_n_680, A2 => gl_ram_n_697, ZN => gl_ram_n_709);
  gl_ram_g55965 : NR2XD2BWP7T port map(A1 => gl_ram_n_691, A2 => gl_ram_n_674, ZN => gl_ram_n_707);
  gl_ram_g55966 : NR2XD2BWP7T port map(A1 => gl_ram_n_688, A2 => gl_ram_n_686, ZN => gl_ram_n_706);
  gl_ram_g55967 : NR2XD3BWP7T port map(A1 => gl_ram_n_685, A2 => gl_ram_n_681, ZN => gl_ram_n_705);
  gl_ram_g55968 : NR2XD3BWP7T port map(A1 => gl_ram_n_690, A2 => gl_ram_n_672, ZN => gl_ram_n_704);
  gl_ram_g55969 : NR2XD3BWP7T port map(A1 => gl_ram_n_678, A2 => gl_ram_n_684, ZN => gl_ram_n_703);
  gl_ram_g55970 : NR2XD2BWP7T port map(A1 => gl_ram_n_689, A2 => gl_ram_n_683, ZN => gl_ram_n_702);
  gl_ram_g55971 : ND2D6BWP7T port map(A1 => gl_ram_n_671, A2 => gl_ram_n_11, ZN => gl_ram_n_701);
  gl_ram_g55974 : MOAI22D0BWP7T port map(A1 => gl_ram_n_664, A2 => FE_PHN528_sig_logic_y_3, B1 => gl_ram_n_664, B2 => FE_PHN516_sig_logic_y_3, ZN => gl_ram_n_698);
  gl_ram_g55975 : AOI21D2BWP7T port map(A1 => gl_ram_n_630, A2 => gl_ram_n_651, B => gl_ram_n_97, ZN => gl_ram_n_697);
  gl_ram_g55977 : INR2D0BWP7T port map(A1 => gl_ram_n_1310, B1 => gl_ram_n_664, ZN => gl_ram_n_695);
  gl_ram_g55982 : AOI21D2BWP7T port map(A1 => gl_ram_n_584, A2 => gl_ram_n_583, B => gl_ram_n_107, ZN => gl_ram_n_690);
  gl_ram_g55983 : AOI21D2BWP7T port map(A1 => gl_ram_n_648, A2 => gl_ram_n_649, B => gl_ram_n_99, ZN => gl_ram_n_689);
  gl_ram_g56002 : AOI21D2BWP7T port map(A1 => gl_ram_n_635, A2 => gl_ram_n_634, B => gl_ram_n_108, ZN => gl_ram_n_676);
  gl_ram_g56003 : AOI21D2BWP7T port map(A1 => gl_ram_n_619, A2 => gl_ram_n_618, B => gl_ram_n_98, ZN => gl_ram_n_675);
  gl_ram_g56004 : AOI21D2BWP7T port map(A1 => gl_ram_n_609, A2 => gl_ram_n_608, B => gl_ram_n_108, ZN => gl_ram_n_674);
  gl_ram_g56006 : AOI21D2BWP7T port map(A1 => gl_ram_n_586, A2 => gl_ram_n_585, B => gl_ram_n_108, ZN => gl_ram_n_672);
  gl_ram_g56019 : MOAI22D0BWP7T port map(A1 => gl_ram_n_611, A2 => gl_ram_n_36, B1 => gl_ram_n_611, B2 => gl_ram_n_36, ZN => gl_ram_n_679);
  gl_ram_g56020 : FA1D0BWP7T port map(A => gl_ram_y_grid(1), B => gl_ram_x_grid(2), CI => gl_ram_n_406, CO => gl_ram_n_662, S => gl_ram_n_663);
  gl_ram_g56021 : HA1D0BWP7T port map(A => FE_PHN530_sig_logic_y_2, B => gl_ram_n_23, CO => gl_ram_n_664, S => gl_ram_n_661);
  gl_ram_g56022 : NR2D2BWP7T port map(A1 => gl_ram_n_577, A2 => gl_ram_n_565, ZN => gl_ram_n_660);
  gl_ram_g56023 : NR2D2BWP7T port map(A1 => gl_ram_n_578, A2 => gl_ram_n_567, ZN => gl_ram_n_659);
  gl_ram_g56024 : NR2XD1BWP7T port map(A1 => gl_ram_n_576, A2 => gl_ram_n_564, ZN => gl_ram_n_658);
  gl_ram_g56026 : ND2D3BWP7T port map(A1 => gl_ram_n_591, A2 => gl_ram_n_613, ZN => gl_ram_n_657);
  gl_ram_g56030 : FA1D0BWP7T port map(A => gl_ram_x_grid(4), B => gl_ram_y_grid(1), CI => gl_ram_y_grid(3), CO => gl_ram_n_652, S => gl_ram_n_653);
  gl_ram_g56031 : NR2XD2BWP7T port map(A1 => gl_ram_n_1483, A2 => gl_ram_n_510, ZN => gl_ram_n_651);
  gl_ram_g56032 : NR2XD2BWP7T port map(A1 => gl_ram_n_1454, A2 => gl_ram_n_548, ZN => gl_ram_n_650);
  gl_ram_g56033 : NR2XD2BWP7T port map(A1 => gl_ram_n_1455, A2 => gl_ram_n_547, ZN => gl_ram_n_649);
  gl_ram_g56034 : NR2XD2BWP7T port map(A1 => gl_ram_n_1456, A2 => gl_ram_n_545, ZN => gl_ram_n_648);
  gl_ram_g56035 : NR2XD2BWP7T port map(A1 => gl_ram_n_1457, A2 => gl_ram_n_543, ZN => gl_ram_n_647);
  gl_ram_g56036 : NR2XD2BWP7T port map(A1 => gl_ram_n_1458, A2 => gl_ram_n_541, ZN => gl_ram_n_646);
  gl_ram_g56037 : NR2XD2BWP7T port map(A1 => gl_ram_n_1460, A2 => gl_ram_n_1459, ZN => gl_ram_n_645);
  gl_ram_g56038 : NR2XD2BWP7T port map(A1 => gl_ram_n_1461, A2 => gl_ram_n_1462, ZN => gl_ram_n_644);
  gl_ram_g56039 : NR2XD2BWP7T port map(A1 => gl_ram_n_1464, A2 => gl_ram_n_1463, ZN => gl_ram_n_643);
  gl_ram_g56040 : NR2XD2BWP7T port map(A1 => gl_ram_n_1466, A2 => gl_ram_n_1465, ZN => gl_ram_n_642);
  gl_ram_g56041 : NR2XD2BWP7T port map(A1 => gl_ram_n_1467, A2 => gl_ram_n_1551, ZN => gl_ram_n_641);
  gl_ram_g56042 : NR2XD2BWP7T port map(A1 => gl_ram_n_1469, A2 => gl_ram_n_1468, ZN => gl_ram_n_640);
  gl_ram_g56043 : NR2XD2BWP7T port map(A1 => gl_ram_n_526, A2 => gl_ram_n_1470, ZN => gl_ram_n_639);
  gl_ram_g56044 : NR2XD2BWP7T port map(A1 => gl_ram_n_1472, A2 => gl_ram_n_1471, ZN => gl_ram_n_638);
  gl_ram_g56045 : NR2D3BWP7T port map(A1 => gl_ram_n_1474, A2 => gl_ram_n_1473, ZN => gl_ram_n_637);
  gl_ram_g56046 : NR2D3BWP7T port map(A1 => gl_ram_n_1476, A2 => gl_ram_n_1475, ZN => gl_ram_n_636);
  gl_ram_g56047 : NR2XD3BWP7T port map(A1 => gl_ram_n_1477, A2 => gl_ram_n_518, ZN => gl_ram_n_635);
  gl_ram_g56048 : NR2XD3BWP7T port map(A1 => gl_ram_n_1478, A2 => gl_ram_n_517, ZN => gl_ram_n_634);
  gl_ram_g56049 : NR2XD3BWP7T port map(A1 => gl_ram_n_1479, A2 => gl_ram_n_1480, ZN => gl_ram_n_633);
  gl_ram_g56050 : NR2XD2BWP7T port map(A1 => gl_ram_n_1482, A2 => gl_ram_n_1481, ZN => gl_ram_n_632);
  gl_ram_g56051 : NR2XD3BWP7T port map(A1 => gl_ram_n_1453, A2 => gl_ram_n_550, ZN => gl_ram_n_631);
  gl_ram_g56052 : NR2XD2BWP7T port map(A1 => gl_ram_n_1484, A2 => gl_ram_n_508, ZN => gl_ram_n_630);
  gl_ram_g56053 : NR2XD2BWP7T port map(A1 => gl_ram_n_1485, A2 => gl_ram_n_507, ZN => gl_ram_n_629);
  gl_ram_g56054 : NR2XD2BWP7T port map(A1 => gl_ram_n_1486, A2 => gl_ram_n_1487, ZN => gl_ram_n_628);
  gl_ram_g56055 : NR2XD2BWP7T port map(A1 => gl_ram_n_1488, A2 => gl_ram_n_503, ZN => gl_ram_n_627);
  gl_ram_g56056 : NR2XD2BWP7T port map(A1 => gl_ram_n_1489, A2 => gl_ram_n_500, ZN => gl_ram_n_626);
  gl_ram_g56057 : NR2D4BWP7T port map(A1 => gl_ram_n_498, A2 => gl_ram_n_499, ZN => gl_ram_n_625);
  gl_ram_g56058 : NR2XD2BWP7T port map(A1 => gl_ram_n_496, A2 => gl_ram_n_1490, ZN => gl_ram_n_624);
  gl_ram_g56059 : NR2XD2BWP7T port map(A1 => gl_ram_n_1452, A2 => gl_ram_n_495, ZN => gl_ram_n_623);
  gl_ram_g56060 : NR2D4BWP7T port map(A1 => gl_ram_n_1494, A2 => gl_ram_n_570, ZN => gl_ram_n_622);
  gl_ram_g56061 : NR2XD2BWP7T port map(A1 => gl_ram_n_1517, A2 => gl_ram_n_571, ZN => gl_ram_n_621);
  gl_ram_g56062 : NR2XD2BWP7T port map(A1 => gl_ram_n_492, A2 => gl_ram_n_1492, ZN => gl_ram_n_620);
  gl_ram_g56063 : NR2XD2BWP7T port map(A1 => gl_ram_n_1496, A2 => gl_ram_n_1497, ZN => gl_ram_n_619);
  gl_ram_g56064 : NR2XD2BWP7T port map(A1 => gl_ram_n_1495, A2 => gl_ram_n_1493, ZN => gl_ram_n_618);
  gl_ram_g56065 : NR2D3BWP7T port map(A1 => gl_ram_n_1498, A2 => gl_ram_n_485, ZN => gl_ram_n_617);
  gl_ram_g56066 : NR2XD2BWP7T port map(A1 => gl_ram_n_1552, A2 => gl_ram_n_484, ZN => gl_ram_n_616);
  gl_ram_g56067 : NR2D3BWP7T port map(A1 => gl_ram_n_482, A2 => gl_ram_n_481, ZN => gl_ram_n_615);
  gl_ram_g56068 : NR2D4BWP7T port map(A1 => gl_ram_n_1501, A2 => gl_ram_n_1499, ZN => gl_ram_n_614);
  gl_ram_g56069 : NR2XD2BWP7T port map(A1 => gl_ram_n_1528, A2 => gl_ram_n_1500, ZN => gl_ram_n_613);
  gl_ram_g56071 : NR2XD2BWP7T port map(A1 => gl_ram_n_1532, A2 => gl_ram_n_1533, ZN => gl_ram_n_610);
  gl_ram_g56072 : NR2XD2BWP7T port map(A1 => gl_ram_n_1507, A2 => gl_ram_n_472, ZN => gl_ram_n_609);
  gl_ram_g56073 : NR2XD2BWP7T port map(A1 => gl_ram_n_467, A2 => gl_ram_n_471, ZN => gl_ram_n_608);
  gl_ram_g56074 : NR2XD2BWP7T port map(A1 => gl_ram_n_1508, A2 => gl_ram_n_1509, ZN => gl_ram_n_607);
  gl_ram_g56075 : NR2XD2BWP7T port map(A1 => gl_ram_n_1510, A2 => gl_ram_n_463, ZN => gl_ram_n_606);
  gl_ram_g56076 : NR2XD2BWP7T port map(A1 => gl_ram_n_1511, A2 => gl_ram_n_459, ZN => gl_ram_n_605);
  gl_ram_g56077 : NR2XD2BWP7T port map(A1 => gl_ram_n_1515, A2 => gl_ram_n_1516, ZN => gl_ram_n_604);
  gl_ram_g56078 : NR2XD2BWP7T port map(A1 => gl_ram_n_457, A2 => gl_ram_n_458, ZN => gl_ram_n_603);
  gl_ram_g56079 : NR2XD2BWP7T port map(A1 => gl_ram_n_1513, A2 => gl_ram_n_1514, ZN => gl_ram_n_602);
  gl_ram_g56080 : NR2XD2BWP7T port map(A1 => gl_ram_n_450, A2 => gl_ram_n_1491, ZN => gl_ram_n_601);
  gl_ram_g56081 : NR2XD2BWP7T port map(A1 => gl_ram_n_1519, A2 => gl_ram_n_1518, ZN => gl_ram_n_600);
  gl_ram_g56082 : NR2XD2BWP7T port map(A1 => gl_ram_n_1520, A2 => gl_ram_n_451, ZN => gl_ram_n_599);
  gl_ram_g56084 : NR2XD2BWP7T port map(A1 => gl_ram_n_1512, A2 => gl_ram_n_1522, ZN => gl_ram_n_597);
  gl_ram_g56085 : NR2XD2BWP7T port map(A1 => gl_ram_n_1524, A2 => gl_ram_n_1523, ZN => gl_ram_n_596);
  gl_ram_g56086 : NR2XD2BWP7T port map(A1 => gl_ram_n_1506, A2 => gl_ram_n_465, ZN => gl_ram_n_595);
  gl_ram_g56087 : NR2D3BWP7T port map(A1 => gl_ram_n_1505, A2 => gl_ram_n_1525, ZN => gl_ram_n_594);
  gl_ram_g56088 : NR2XD2BWP7T port map(A1 => gl_ram_n_1526, A2 => gl_ram_n_1502, ZN => gl_ram_n_593);
  gl_ram_g56089 : NR2XD2BWP7T port map(A1 => gl_ram_n_1527, A2 => gl_ram_n_439, ZN => gl_ram_n_592);
  gl_ram_g56090 : NR2XD2BWP7T port map(A1 => gl_ram_n_1530, A2 => gl_ram_n_1529, ZN => gl_ram_n_591);
  gl_ram_g56091 : NR2XD2BWP7T port map(A1 => gl_ram_n_1504, A2 => gl_ram_n_1503, ZN => gl_ram_n_590);
  gl_ram_g56092 : NR2XD2BWP7T port map(A1 => gl_ram_n_433, A2 => gl_ram_n_1531, ZN => gl_ram_n_589);
  gl_ram_g56093 : NR2XD3BWP7T port map(A1 => gl_ram_n_1535, A2 => gl_ram_n_1534, ZN => gl_ram_n_588);
  gl_ram_g56094 : NR2XD2BWP7T port map(A1 => gl_ram_n_1537, A2 => gl_ram_n_1536, ZN => gl_ram_n_587);
  gl_ram_g56095 : NR2XD3BWP7T port map(A1 => gl_ram_n_1538, A2 => gl_ram_n_424, ZN => gl_ram_n_586);
  gl_ram_g56096 : NR2XD2BWP7T port map(A1 => gl_ram_n_1539, A2 => gl_ram_n_426, ZN => gl_ram_n_585);
  gl_ram_g56097 : NR2XD3BWP7T port map(A1 => gl_ram_n_1540, A2 => gl_ram_n_1541, ZN => gl_ram_n_584);
  gl_ram_g56098 : NR2XD3BWP7T port map(A1 => gl_ram_n_1543, A2 => gl_ram_n_1542, ZN => gl_ram_n_583);
  gl_ram_g56099 : NR2XD2BWP7T port map(A1 => gl_ram_n_1544, A2 => gl_ram_n_417, ZN => gl_ram_n_582);
  gl_ram_g56100 : NR2XD2BWP7T port map(A1 => gl_ram_n_1545, A2 => gl_ram_n_415, ZN => gl_ram_n_581);
  gl_ram_g56101 : NR2XD2BWP7T port map(A1 => gl_ram_n_1548, A2 => gl_ram_n_1547, ZN => gl_ram_n_580);
  gl_ram_g56102 : NR2XD2BWP7T port map(A1 => gl_ram_n_1546, A2 => gl_ram_n_414, ZN => gl_ram_n_579);
  gl_ram_g56103 : OAI21D2BWP7T port map(A1 => gl_ram_n_14, A2 => gl_ram_n_258, B => gl_ram_n_111, ZN => gl_ram_n_578);
  gl_ram_g56104 : OAI21D2BWP7T port map(A1 => gl_ram_n_20, A2 => gl_ram_n_258, B => gl_ram_n_112, ZN => gl_ram_n_577);
  gl_ram_g56105 : OAI21D2BWP7T port map(A1 => gl_ram_n_15, A2 => gl_ram_n_259, B => gl_ram_n_110, ZN => gl_ram_n_576);
  gl_ram_g56106 : NR2XD1BWP7T port map(A1 => gl_ram_n_3, A2 => gl_ram_n_568, ZN => gl_ram_n_575);
  gl_ram_g56108 : NR2XD2BWP7T port map(A1 => gl_ram_n_2, A2 => gl_ram_n_1450, ZN => gl_ram_n_573);
  gl_ram_g56109 : MOAI22D0BWP7T port map(A1 => gl_ram_n_24, A2 => sig_logic_x(3), B1 => gl_ram_n_24, B2 => sig_logic_x(3), ZN => gl_ram_n_572);
  gl_ram_g56110 : CKXOR2D0BWP7T port map(A1 => gl_ram_y_grid(3), A2 => gl_ram_n_113, Z => gl_ram_n_611);
  gl_ram_g56111 : ND2D2BWP7T port map(A1 => gl_ram_n_285, A2 => gl_ram_n_286, ZN => gl_ram_n_571);
  gl_ram_g56112 : ND2D3BWP7T port map(A1 => gl_ram_n_270, A2 => gl_ram_n_272, ZN => gl_ram_n_570);
  gl_ram_g56115 : AN2D4BWP7T port map(A1 => gl_ram_ram_96(2), A2 => gl_ram_n_6, Z => gl_ram_n_568);
  gl_ram_g56116 : AN2D2BWP7T port map(A1 => gl_ram_ram_99(2), A2 => gl_ram_n_5, Z => gl_ram_n_567);
  gl_ram_g56119 : NR2D3BWP7T port map(A1 => gl_ram_n_1440, A2 => gl_ram_n_259, ZN => gl_ram_n_565);
  gl_ram_g56121 : AN2XD1BWP7T port map(A1 => gl_ram_ram_96(1), A2 => gl_ram_n_6, Z => gl_ram_n_564);
  gl_ram_g56123 : NR2D1BWP7T port map(A1 => gl_ram_n_408, A2 => gl_ram_n_96, ZN => gl_ram_n_563);
  gl_ram_g56124 : OR2D1BWP7T port map(A1 => gl_ram_n_409, A2 => gl_ram_n_96, Z => gl_ram_n_562);
  gl_ram_g56125 : OR2D1BWP7T port map(A1 => gl_ram_n_256, A2 => gl_ram_n_96, Z => gl_ram_n_561);
  gl_ram_g56126 : OR2D1BWP7T port map(A1 => gl_ram_n_408, A2 => gl_ram_n_98, Z => gl_ram_n_560);
  gl_ram_g56127 : NR2XD0BWP7T port map(A1 => gl_ram_n_408, A2 => gl_ram_n_99, ZN => gl_ram_n_559);
  gl_ram_g56128 : OR2D1BWP7T port map(A1 => gl_ram_n_408, A2 => gl_ram_n_97, Z => gl_ram_n_558);
  gl_ram_g56129 : OR2D1BWP7T port map(A1 => gl_ram_n_409, A2 => gl_ram_n_98, Z => gl_ram_n_557);
  gl_ram_g56130 : OR2D1BWP7T port map(A1 => gl_ram_n_409, A2 => gl_ram_n_99, Z => gl_ram_n_556);
  gl_ram_g56131 : NR2D1BWP7T port map(A1 => gl_ram_n_256, A2 => gl_ram_n_98, ZN => gl_ram_n_555);
  gl_ram_g56132 : OR2D1BWP7T port map(A1 => gl_ram_n_409, A2 => gl_ram_n_97, Z => gl_ram_n_554);
  gl_ram_g56133 : NR2XD0BWP7T port map(A1 => gl_ram_n_256, A2 => gl_ram_n_99, ZN => gl_ram_n_553);
  gl_ram_g56134 : OR2D1BWP7T port map(A1 => gl_ram_n_256, A2 => gl_ram_n_97, Z => gl_ram_n_552);
  gl_ram_g56136 : ND2D3BWP7T port map(A1 => gl_ram_n_399, A2 => gl_ram_n_400, ZN => gl_ram_n_550);
  gl_ram_g56138 : ND2D2BWP7T port map(A1 => gl_ram_n_396, A2 => gl_ram_n_395, ZN => gl_ram_n_548);
  gl_ram_g56139 : ND2D2BWP7T port map(A1 => gl_ram_n_393, A2 => gl_ram_n_394, ZN => gl_ram_n_547);
  gl_ram_g56141 : ND2D2BWP7T port map(A1 => gl_ram_n_389, A2 => gl_ram_n_390, ZN => gl_ram_n_545);
  gl_ram_g56145 : ND2D2BWP7T port map(A1 => gl_ram_n_379, A2 => gl_ram_n_380, ZN => gl_ram_n_541);
  gl_ram_g56160 : IOA21D2BWP7T port map(A1 => gl_ram_ram_80(2), A2 => gl_ram_n_89, B => gl_ram_n_348, ZN => gl_ram_n_526);
  gl_ram_g56168 : ND2D3BWP7T port map(A1 => gl_ram_n_332, A2 => gl_ram_n_333, ZN => gl_ram_n_518);
  gl_ram_g56169 : ND2D3BWP7T port map(A1 => gl_ram_n_330, A2 => gl_ram_n_331, ZN => gl_ram_n_517);
  gl_ram_g56179 : ND2D2BWP7T port map(A1 => gl_ram_n_309, A2 => gl_ram_n_310, ZN => gl_ram_n_507);
  gl_ram_g56183 : ND2D3BWP7T port map(A1 => gl_ram_n_301, A2 => gl_ram_n_300, ZN => gl_ram_n_503);
  gl_ram_g56186 : ND2D3BWP7T port map(A1 => gl_ram_n_164, A2 => gl_ram_n_296, ZN => gl_ram_n_500);
  gl_ram_g56187 : ND2D2BWP7T port map(A1 => gl_ram_n_297, A2 => gl_ram_n_293, ZN => gl_ram_n_499);
  gl_ram_g56188 : ND2D3BWP7T port map(A1 => gl_ram_n_291, A2 => gl_ram_n_288, ZN => gl_ram_n_498);
  gl_ram_g56190 : ND2D2BWP7T port map(A1 => gl_ram_n_294, A2 => gl_ram_n_156, ZN => gl_ram_n_496);
  gl_ram_g56191 : ND2D3BWP7T port map(A1 => gl_ram_n_290, A2 => gl_ram_n_289, ZN => gl_ram_n_495);
  gl_ram_g56197 : ND2D2BWP7T port map(A1 => gl_ram_n_281, A2 => gl_ram_n_282, ZN => gl_ram_n_492);
  gl_ram_g56204 : ND2D3BWP7T port map(A1 => gl_ram_n_264, A2 => gl_ram_n_263, ZN => gl_ram_n_485);
  gl_ram_g56205 : ND2D3BWP7T port map(A1 => gl_ram_n_260, A2 => gl_ram_n_261, ZN => gl_ram_n_484);
  gl_ram_g56207 : ND2D2BWP7T port map(A1 => gl_ram_n_254, A2 => gl_ram_n_403, ZN => gl_ram_n_482);
  gl_ram_g56208 : ND2D2BWP7T port map(A1 => gl_ram_n_252, A2 => gl_ram_n_253, ZN => gl_ram_n_481);
  gl_ram_g56214 : ND2D2BWP7T port map(A1 => gl_ram_n_241, A2 => gl_ram_n_242, ZN => gl_ram_n_475);
  gl_ram_g56217 : ND2D2BWP7T port map(A1 => gl_ram_n_228, A2 => gl_ram_n_227, ZN => gl_ram_n_472);
  gl_ram_g56218 : ND2D2BWP7T port map(A1 => gl_ram_n_226, A2 => gl_ram_n_224, ZN => gl_ram_n_471);
  gl_ram_g56222 : ND2D2BWP7T port map(A1 => gl_ram_n_222, A2 => gl_ram_n_221, ZN => gl_ram_n_467);
  gl_ram_g56224 : ND2D2BWP7T port map(A1 => gl_ram_n_225, A2 => gl_ram_n_231, ZN => gl_ram_n_465);
  gl_ram_g56226 : ND2D2BWP7T port map(A1 => gl_ram_n_215, A2 => gl_ram_n_214, ZN => gl_ram_n_463);
  gl_ram_g56231 : ND2D3BWP7T port map(A1 => gl_ram_n_204, A2 => gl_ram_n_203, ZN => gl_ram_n_458);
  gl_ram_g56232 : ND2D2BWP7T port map(A1 => gl_ram_n_201, A2 => gl_ram_n_202, ZN => gl_ram_n_457);
  gl_ram_g56238 : ND2D2BWP7T port map(A1 => gl_ram_n_255, A2 => gl_ram_n_189, ZN => gl_ram_n_451);
  gl_ram_g56239 : ND2D2BWP7T port map(A1 => gl_ram_n_186, A2 => gl_ram_n_187, ZN => gl_ram_n_450);
  gl_ram_g56250 : ND2D2BWP7T port map(A1 => gl_ram_n_246, A2 => gl_ram_n_169, ZN => gl_ram_n_439);
  gl_ram_g56256 : IOA21D2BWP7T port map(A1 => gl_ram_ram_81(1), A2 => gl_ram_n_88, B => gl_ram_n_312, ZN => gl_ram_n_433);
  gl_ram_g56265 : ND2D4BWP7T port map(A1 => gl_ram_n_145, A2 => gl_ram_n_143, ZN => gl_ram_n_424);
  gl_ram_g56272 : ND2D3BWP7T port map(A1 => gl_ram_n_128, A2 => gl_ram_n_126, ZN => gl_ram_n_417);
  gl_ram_g56274 : ND2D3BWP7T port map(A1 => gl_ram_n_125, A2 => gl_ram_n_124, ZN => gl_ram_n_415);
  gl_ram_g56275 : ND2D2BWP7T port map(A1 => gl_ram_n_121, A2 => gl_ram_n_120, ZN => gl_ram_n_414);
  gl_ram_g56279 : MOAI22D0BWP7T port map(A1 => gl_ram_n_36, A2 => gl_ram_y_grid(2), B1 => gl_ram_n_36, B2 => gl_ram_y_grid(2), ZN => gl_ram_n_410);
  gl_ram_g56280 : HA1D0BWP7T port map(A => gl_ram_x_grid(1), B => gl_ram_y_grid(0), CO => gl_ram_n_406, S => gl_ram_n_407);
  gl_ram_g56281 : HA1D0BWP7T port map(A => gl_ram_x_grid(3), B => gl_ram_y_grid(0), CO => gl_ram_n_404, S => gl_ram_n_405);
  gl_ram_g56282 : ND2D2BWP7T port map(A1 => gl_ram_ram_87(0), A2 => gl_ram_n_92, ZN => gl_ram_n_403);
  gl_ram_g56284 : CKND2D2BWP7T port map(A1 => gl_ram_ram_15(1), A2 => gl_ram_n_92, ZN => gl_ram_n_401);
  gl_ram_g56285 : CKND2D2BWP7T port map(A1 => gl_ram_ram_14(1), A2 => gl_ram_n_93, ZN => gl_ram_n_400);
  gl_ram_g56286 : CKND2D2BWP7T port map(A1 => gl_ram_ram_12(1), A2 => gl_ram_n_91, ZN => gl_ram_n_399);
  gl_ram_g56287 : ND2D2BWP7T port map(A1 => gl_ram_ram_10(1), A2 => gl_ram_n_86, ZN => gl_ram_n_398);
  gl_ram_g56289 : CKND2D2BWP7T port map(A1 => gl_ram_ram_11(1), A2 => gl_ram_n_87, ZN => gl_ram_n_396);
  gl_ram_g56290 : CKND2D2BWP7T port map(A1 => gl_ram_ram_8(1), A2 => gl_ram_n_89, ZN => gl_ram_n_395);
  gl_ram_g56291 : ND2D2BWP7T port map(A1 => gl_ram_ram_21(1), A2 => gl_ram_n_90, ZN => gl_ram_n_394);
  gl_ram_g56292 : ND2D2BWP7T port map(A1 => gl_ram_ram_23(1), A2 => gl_ram_n_92, ZN => gl_ram_n_393);
  gl_ram_g56294 : ND2D2BWP7T port map(A1 => gl_ram_ram_20(1), A2 => gl_ram_n_91, ZN => gl_ram_n_391);
  gl_ram_g56295 : CKND2D2BWP7T port map(A1 => gl_ram_ram_18(1), A2 => gl_ram_n_86, ZN => gl_ram_n_390);
  gl_ram_g56296 : CKND2D2BWP7T port map(A1 => gl_ram_ram_17(1), A2 => gl_ram_n_88, ZN => gl_ram_n_389);
  gl_ram_g56297 : CKND2D2BWP7T port map(A1 => gl_ram_ram_19(1), A2 => gl_ram_n_87, ZN => gl_ram_n_388);
  gl_ram_g56298 : ND2D2BWP7T port map(A1 => gl_ram_ram_3(1), A2 => gl_ram_n_87, ZN => gl_ram_n_387);
  gl_ram_g56304 : ND2D2BWP7T port map(A1 => gl_ram_ram_52(1), A2 => gl_ram_n_91, ZN => gl_ram_n_381);
  gl_ram_g56305 : ND2D2BWP7T port map(A1 => gl_ram_ram_49(1), A2 => gl_ram_n_88, ZN => gl_ram_n_380);
  gl_ram_g56307 : ND2D2BWP7T port map(A1 => gl_ram_ram_51(1), A2 => gl_ram_n_87, ZN => gl_ram_n_378);
  gl_ram_g56312 : ND2D2BWP7T port map(A1 => gl_ram_ram_4(1), A2 => gl_ram_n_91, ZN => gl_ram_n_373);
  gl_ram_g56314 : ND2D2BWP7T port map(A1 => gl_ram_ram_2(1), A2 => gl_ram_n_86, ZN => gl_ram_n_371);
  gl_ram_g56319 : CKND2D2BWP7T port map(A1 => gl_ram_ram_79(2), A2 => gl_ram_n_92, ZN => gl_ram_n_366);
  gl_ram_g56323 : CKND2D2BWP7T port map(A1 => gl_ram_ram_76(2), A2 => gl_ram_n_91, ZN => gl_ram_n_362);
  gl_ram_g56324 : ND2D2BWP7T port map(A1 => gl_ram_ram_75(2), A2 => gl_ram_n_87, ZN => gl_ram_n_361);
  gl_ram_g56325 : ND2D2BWP7T port map(A1 => gl_ram_ram_36(2), A2 => gl_ram_n_91, ZN => gl_ram_n_360);
  gl_ram_g56326 : CKND2D2BWP7T port map(A1 => gl_ram_ram_71(2), A2 => gl_ram_n_92, ZN => gl_ram_n_359);
  gl_ram_g56328 : ND2D2BWP7T port map(A1 => gl_ram_ram_68(2), A2 => gl_ram_n_91, ZN => gl_ram_n_357);
  gl_ram_g56331 : ND2D2BWP7T port map(A1 => gl_ram_ram_66(2), A2 => gl_ram_n_86, ZN => gl_ram_n_354);
  gl_ram_g56332 : CKND2D2BWP7T port map(A1 => gl_ram_ram_67(2), A2 => gl_ram_n_87, ZN => gl_ram_n_353);
  gl_ram_g56334 : CKND2D2BWP7T port map(A1 => gl_ram_ram_87(2), A2 => gl_ram_n_92, ZN => gl_ram_n_351);
  gl_ram_g56335 : ND2D2BWP7T port map(A1 => gl_ram_ram_24(2), A2 => gl_ram_n_89, ZN => gl_ram_n_350);
  gl_ram_g56337 : ND2D2BWP7T port map(A1 => gl_ram_ram_83(2), A2 => gl_ram_n_87, ZN => gl_ram_n_348);
  gl_ram_g56339 : ND2D2BWP7T port map(A1 => gl_ram_ram_84(2), A2 => gl_ram_n_91, ZN => gl_ram_n_346);
  gl_ram_g56340 : ND2D2BWP7T port map(A1 => gl_ram_ram_82(2), A2 => gl_ram_n_86, ZN => gl_ram_n_345);
  gl_ram_g56342 : ND2D2BWP7T port map(A1 => gl_ram_ram_95(2), A2 => gl_ram_n_92, ZN => gl_ram_n_343);
  gl_ram_g56345 : ND2D1BWP7T port map(A1 => gl_ram_ram_92(2), A2 => gl_ram_n_91, ZN => gl_ram_n_340);
  gl_ram_g56346 : ND2D2BWP7T port map(A1 => gl_ram_ram_90(2), A2 => gl_ram_n_86, ZN => gl_ram_n_339);
  gl_ram_g56349 : ND2D2BWP7T port map(A1 => gl_ram_ram_91(2), A2 => gl_ram_n_87, ZN => gl_ram_n_336);
  gl_ram_g56350 : ND2D2BWP7T port map(A1 => gl_ram_ram_63(2), A2 => gl_ram_n_92, ZN => gl_ram_n_335);
  gl_ram_g56352 : ND2D2BWP7T port map(A1 => gl_ram_ram_62(2), A2 => gl_ram_n_93, ZN => gl_ram_n_333);
  gl_ram_g56353 : ND2D2BWP7T port map(A1 => gl_ram_ram_60(2), A2 => gl_ram_n_91, ZN => gl_ram_n_332);
  gl_ram_g56354 : ND2D2BWP7T port map(A1 => gl_ram_ram_58(2), A2 => gl_ram_n_86, ZN => gl_ram_n_331);
  gl_ram_g56355 : CKND2D3BWP7T port map(A1 => gl_ram_ram_57(2), A2 => gl_ram_n_88, ZN => gl_ram_n_330);
  gl_ram_g56359 : ND2D2BWP7T port map(A1 => gl_ram_ram_47(2), A2 => gl_ram_n_92, ZN => gl_ram_n_326);
  gl_ram_g56363 : ND2D2BWP7T port map(A1 => gl_ram_ram_41(2), A2 => gl_ram_n_88, ZN => gl_ram_n_322);
  gl_ram_g56369 : ND2D2BWP7T port map(A1 => gl_ram_ram_28(2), A2 => gl_ram_n_91, ZN => gl_ram_n_316);
  gl_ram_g56370 : ND2D2BWP7T port map(A1 => gl_ram_ram_26(2), A2 => gl_ram_n_86, ZN => gl_ram_n_315);
  gl_ram_g56373 : ND2D2BWP7T port map(A1 => gl_ram_ram_82(1), A2 => gl_ram_n_86, ZN => gl_ram_n_312);
  gl_ram_g56374 : ND2D2BWP7T port map(A1 => gl_ram_ram_19(2), A2 => gl_ram_n_87, ZN => gl_ram_n_311);
  gl_ram_g56375 : ND2D2BWP7T port map(A1 => gl_ram_ram_39(2), A2 => gl_ram_n_92, ZN => gl_ram_n_310);
  gl_ram_g56376 : ND2D2BWP7T port map(A1 => gl_ram_ram_37(2), A2 => gl_ram_n_90, ZN => gl_ram_n_309);
  gl_ram_g56378 : ND2D2BWP7T port map(A1 => gl_ram_ram_34(2), A2 => gl_ram_n_86, ZN => gl_ram_n_307);
  gl_ram_g56380 : ND2D2BWP7T port map(A1 => gl_ram_ram_35(2), A2 => gl_ram_n_87, ZN => gl_ram_n_305);
  gl_ram_g56381 : ND2D2BWP7T port map(A1 => gl_ram_ram_67(0), A2 => gl_ram_n_87, ZN => gl_ram_n_304);
  gl_ram_g56382 : ND2D2BWP7T port map(A1 => gl_ram_ram_15(2), A2 => gl_ram_n_92, ZN => gl_ram_n_303);
  gl_ram_g56384 : ND2D2BWP7T port map(A1 => gl_ram_ram_12(2), A2 => gl_ram_n_91, ZN => gl_ram_n_301);
  gl_ram_g56385 : ND2D2BWP7T port map(A1 => gl_ram_ram_14(2), A2 => gl_ram_n_93, ZN => gl_ram_n_300);
  gl_ram_g56386 : ND2D2BWP7T port map(A1 => gl_ram_ram_10(2), A2 => gl_ram_n_86, ZN => gl_ram_n_299);
  gl_ram_g56388 : ND2D2BWP7T port map(A1 => gl_ram_ram_79(0), A2 => gl_ram_n_92, ZN => gl_ram_n_297);
  gl_ram_g56389 : ND2D2BWP7T port map(A1 => gl_ram_ram_8(2), A2 => gl_ram_n_89, ZN => gl_ram_n_296);
  gl_ram_g56391 : ND2D2BWP7T port map(A1 => gl_ram_ram_23(2), A2 => gl_ram_n_92, ZN => gl_ram_n_294);
  gl_ram_g56392 : CKND2D2BWP7T port map(A1 => gl_ram_ram_77(0), A2 => gl_ram_n_90, ZN => gl_ram_n_293);
  gl_ram_g56393 : ND2D2BWP7T port map(A1 => gl_ram_ram_20(2), A2 => gl_ram_n_91, ZN => gl_ram_n_292);
  gl_ram_g56394 : ND2D2BWP7T port map(A1 => gl_ram_ram_78(0), A2 => gl_ram_n_93, ZN => gl_ram_n_291);
  gl_ram_g56395 : ND2D2BWP7T port map(A1 => gl_ram_ram_17(2), A2 => gl_ram_n_88, ZN => gl_ram_n_290);
  gl_ram_g56396 : ND2D2BWP7T port map(A1 => gl_ram_ram_18(2), A2 => gl_ram_n_86, ZN => gl_ram_n_289);
  gl_ram_g56397 : ND2D2BWP7T port map(A1 => gl_ram_ram_76(0), A2 => gl_ram_n_91, ZN => gl_ram_n_288);
  gl_ram_g56399 : ND2D2BWP7T port map(A1 => gl_ram_ram_55(2), A2 => gl_ram_n_92, ZN => gl_ram_n_286);
  gl_ram_g56400 : ND2D2BWP7T port map(A1 => gl_ram_ram_53(2), A2 => gl_ram_n_90, ZN => gl_ram_n_285);
  gl_ram_g56406 : ND2D2BWP7T port map(A1 => gl_ram_ram_51(2), A2 => gl_ram_n_87, ZN => gl_ram_n_279);
  gl_ram_g56408 : ND2D2BWP7T port map(A1 => gl_ram_ram_75(0), A2 => gl_ram_n_87, ZN => gl_ram_n_277);
  gl_ram_g56409 : ND2D2BWP7T port map(A1 => gl_ram_ram_7(2), A2 => gl_ram_n_92, ZN => gl_ram_n_276);
  gl_ram_g56411 : ND2D2BWP7T port map(A1 => gl_ram_ram_4(2), A2 => gl_ram_n_91, ZN => gl_ram_n_274);
  gl_ram_g56412 : ND2D2BWP7T port map(A1 => gl_ram_ram_2(2), A2 => gl_ram_n_86, ZN => gl_ram_n_273);
  gl_ram_g56413 : ND2D3BWP7T port map(A1 => gl_ram_ram_74(0), A2 => gl_ram_n_86, ZN => gl_ram_n_272);
  gl_ram_g56414 : ND2D2BWP7T port map(A1 => gl_ram_ram_3(2), A2 => gl_ram_n_87, ZN => gl_ram_n_271);
  gl_ram_g56415 : ND2D3BWP7T port map(A1 => gl_ram_ram_73(0), A2 => gl_ram_n_88, ZN => gl_ram_n_270);
  gl_ram_g56416 : ND2D2BWP7T port map(A1 => gl_ram_ram_76(1), A2 => gl_ram_n_91, ZN => gl_ram_n_269);
  gl_ram_g56418 : CKND2D2BWP7T port map(A1 => gl_ram_ram_71(1), A2 => gl_ram_n_92, ZN => gl_ram_n_267);
  gl_ram_g56420 : CKND2D2BWP7T port map(A1 => gl_ram_ram_71(0), A2 => gl_ram_n_92, ZN => gl_ram_n_265);
  gl_ram_g56421 : CKND2D2BWP7T port map(A1 => gl_ram_ram_70(0), A2 => gl_ram_n_93, ZN => gl_ram_n_264);
  gl_ram_g56422 : CKND2D3BWP7T port map(A1 => gl_ram_ram_68(0), A2 => gl_ram_n_91, ZN => gl_ram_n_263);
  gl_ram_g56424 : ND2D3BWP7T port map(A1 => gl_ram_ram_66(0), A2 => gl_ram_n_86, ZN => gl_ram_n_261);
  gl_ram_g56425 : ND2D3BWP7T port map(A1 => gl_ram_ram_65(0), A2 => gl_ram_n_88, ZN => gl_ram_n_260);
  gl_ram_g56427 : AN2D2BWP7T port map(A1 => gl_ram_n_106, A2 => gl_ram_n_112, Z => gl_ram_n_409);
  gl_ram_g56428 : AN2D1BWP7T port map(A1 => gl_ram_n_106, A2 => gl_ram_n_111, Z => gl_ram_n_408);
  gl_ram_g56430 : CKND2D2BWP7T port map(A1 => gl_ram_ram_21(0), A2 => gl_ram_n_90, ZN => gl_ram_n_255);
  gl_ram_g56431 : ND2D2BWP7T port map(A1 => gl_ram_ram_85(0), A2 => gl_ram_n_90, ZN => gl_ram_n_254);
  gl_ram_g56432 : CKND2D3BWP7T port map(A1 => gl_ram_ram_86(0), A2 => gl_ram_n_93, ZN => gl_ram_n_253);
  gl_ram_g56433 : ND2D2BWP7T port map(A1 => gl_ram_ram_84(0), A2 => gl_ram_n_91, ZN => gl_ram_n_252);
  gl_ram_g56434 : CKND2D3BWP7T port map(A1 => gl_ram_ram_82(0), A2 => gl_ram_n_86, ZN => gl_ram_n_251);
  gl_ram_g56436 : ND2D2BWP7T port map(A1 => gl_ram_ram_83(0), A2 => gl_ram_n_87, ZN => gl_ram_n_249);
  gl_ram_g56439 : CKND2D2BWP7T port map(A1 => gl_ram_ram_73(1), A2 => gl_ram_n_88, ZN => gl_ram_n_246);
  gl_ram_g56440 : ND2D2BWP7T port map(A1 => gl_ram_ram_66(1), A2 => gl_ram_n_86, ZN => gl_ram_n_245);
  gl_ram_g56442 : ND2D2BWP7T port map(A1 => gl_ram_ram_79(1), A2 => gl_ram_n_92, ZN => gl_ram_n_243);
  gl_ram_g56443 : ND2D2BWP7T port map(A1 => gl_ram_ram_95(0), A2 => gl_ram_n_92, ZN => gl_ram_n_242);
  gl_ram_g56444 : ND2D2BWP7T port map(A1 => gl_ram_ram_93(0), A2 => gl_ram_n_90, ZN => gl_ram_n_241);
  gl_ram_g56445 : ND2D2BWP7T port map(A1 => gl_ram_ram_35(1), A2 => gl_ram_n_87, ZN => gl_ram_n_240);
  gl_ram_g56446 : ND2D2BWP7T port map(A1 => gl_ram_ram_92(0), A2 => gl_ram_n_91, ZN => gl_ram_n_239);
  gl_ram_g56450 : ND2D2BWP7T port map(A1 => gl_ram_ram_91(0), A2 => gl_ram_n_87, ZN => gl_ram_n_235);
  gl_ram_g56453 : ND2D2BWP7T port map(A1 => gl_ram_ram_90(0), A2 => gl_ram_n_86, ZN => gl_ram_n_232);
  gl_ram_g56454 : ND2D2BWP7T port map(A1 => gl_ram_ram_7(0), A2 => gl_ram_n_92, ZN => gl_ram_n_231);
  gl_ram_g56456 : CKND2D2BWP7T port map(A1 => gl_ram_ram_60(0), A2 => gl_ram_n_91, ZN => gl_ram_n_229);
  gl_ram_g56457 : ND2D2BWP7T port map(A1 => gl_ram_ram_63(0), A2 => gl_ram_n_92, ZN => gl_ram_n_228);
  gl_ram_g56458 : CKND2D2BWP7T port map(A1 => gl_ram_ram_61(0), A2 => gl_ram_n_90, ZN => gl_ram_n_227);
  gl_ram_g56459 : CKND2D2BWP7T port map(A1 => gl_ram_ram_58(0), A2 => gl_ram_n_86, ZN => gl_ram_n_226);
  gl_ram_g56460 : ND2D2BWP7T port map(A1 => gl_ram_ram_5(0), A2 => gl_ram_n_90, ZN => gl_ram_n_225);
  gl_ram_g56461 : ND2D2BWP7T port map(A1 => gl_ram_ram_57(0), A2 => gl_ram_n_88, ZN => gl_ram_n_224);
  gl_ram_g56463 : ND2D2BWP7T port map(A1 => gl_ram_ram_59(0), A2 => gl_ram_n_87, ZN => gl_ram_n_222);
  gl_ram_g56464 : ND2D2BWP7T port map(A1 => gl_ram_ram_56(0), A2 => gl_ram_n_89, ZN => gl_ram_n_221);
  gl_ram_g56465 : ND2D2BWP7T port map(A1 => gl_ram_ram_47(0), A2 => gl_ram_n_92, ZN => gl_ram_n_220);
  gl_ram_g56467 : ND2D2BWP7T port map(A1 => gl_ram_ram_44(0), A2 => gl_ram_n_91, ZN => gl_ram_n_218);
  gl_ram_g56471 : ND2D2BWP7T port map(A1 => gl_ram_ram_41(0), A2 => gl_ram_n_88, ZN => gl_ram_n_214);
  gl_ram_g56472 : ND2D2BWP7T port map(A1 => gl_ram_ram_43(0), A2 => gl_ram_n_87, ZN => gl_ram_n_213);
  gl_ram_g56478 : ND2D2BWP7T port map(A1 => gl_ram_ram_28(0), A2 => gl_ram_n_91, ZN => gl_ram_n_207);
  gl_ram_g56480 : ND2D2BWP7T port map(A1 => gl_ram_ram_31(0), A2 => gl_ram_n_92, ZN => gl_ram_n_205);
  gl_ram_g56481 : CKND2D2BWP7T port map(A1 => gl_ram_ram_25(0), A2 => gl_ram_n_88, ZN => gl_ram_n_204);
  gl_ram_g56482 : ND2D2BWP7T port map(A1 => gl_ram_ram_26(0), A2 => gl_ram_n_86, ZN => gl_ram_n_203);
  gl_ram_g56483 : ND2D2BWP7T port map(A1 => gl_ram_ram_24(0), A2 => gl_ram_n_89, ZN => gl_ram_n_202);
  gl_ram_g56484 : ND2D2BWP7T port map(A1 => gl_ram_ram_27(0), A2 => gl_ram_n_87, ZN => gl_ram_n_201);
  gl_ram_g56491 : ND2D2BWP7T port map(A1 => gl_ram_ram_33(0), A2 => gl_ram_n_88, ZN => gl_ram_n_194);
  gl_ram_g56493 : ND2D2BWP7T port map(A1 => gl_ram_ram_18(0), A2 => gl_ram_n_86, ZN => gl_ram_n_192);
  gl_ram_g56494 : ND2D2BWP7T port map(A1 => gl_ram_ram_35(0), A2 => gl_ram_n_87, ZN => gl_ram_n_191);
  gl_ram_g56496 : ND2D2BWP7T port map(A1 => gl_ram_ram_23(0), A2 => gl_ram_n_92, ZN => gl_ram_n_189);
  gl_ram_g56497 : ND2D2BWP7T port map(A1 => gl_ram_ram_15(0), A2 => gl_ram_n_92, ZN => gl_ram_n_188);
  gl_ram_g56498 : ND2D2BWP7T port map(A1 => gl_ram_ram_14(0), A2 => gl_ram_n_93, ZN => gl_ram_n_187);
  gl_ram_g56499 : ND2D2BWP7T port map(A1 => gl_ram_ram_12(0), A2 => gl_ram_n_91, ZN => gl_ram_n_186);
  gl_ram_g56500 : ND2D2BWP7T port map(A1 => gl_ram_ram_10(0), A2 => gl_ram_n_86, ZN => gl_ram_n_185);
  gl_ram_g56502 : ND2D2BWP7T port map(A1 => gl_ram_ram_11(0), A2 => gl_ram_n_87, ZN => gl_ram_n_183);
  gl_ram_g56504 : ND2D2BWP7T port map(A1 => gl_ram_ram_91(1), A2 => gl_ram_n_87, ZN => gl_ram_n_181);
  gl_ram_g56506 : ND2D2BWP7T port map(A1 => gl_ram_ram_20(0), A2 => gl_ram_n_91, ZN => gl_ram_n_179);
  gl_ram_g56507 : ND2D2BWP7T port map(A1 => gl_ram_ram_19(0), A2 => gl_ram_n_87, ZN => gl_ram_n_178);
  gl_ram_g56511 : ND2D2BWP7T port map(A1 => gl_ram_ram_36(0), A2 => gl_ram_n_91, ZN => gl_ram_n_174);
  gl_ram_g56512 : ND2D2BWP7T port map(A1 => gl_ram_ram_2(0), A2 => gl_ram_n_86, ZN => gl_ram_n_173);
  gl_ram_g56514 : ND2D1P5BWP7T port map(A1 => gl_ram_ram_3(0), A2 => gl_ram_n_87, ZN => gl_ram_n_171);
  gl_ram_g56516 : ND2D1BWP7T port map(A1 => gl_ram_ram_74(1), A2 => gl_ram_n_86, ZN => gl_ram_n_169);
  gl_ram_g56517 : ND2D2BWP7T port map(A1 => gl_ram_ram_75(1), A2 => gl_ram_n_87, ZN => gl_ram_n_168);
  gl_ram_g56519 : ND2D2BWP7T port map(A1 => gl_ram_ram_67(1), A2 => gl_ram_n_87, ZN => gl_ram_n_166);
  gl_ram_g56521 : ND2D2BWP7T port map(A1 => gl_ram_ram_11(2), A2 => gl_ram_n_87, ZN => gl_ram_n_164);
  gl_ram_g56522 : ND2D2BWP7T port map(A1 => gl_ram_ram_68(1), A2 => gl_ram_n_91, ZN => gl_ram_n_163);
  gl_ram_g56523 : ND2D2BWP7T port map(A1 => gl_ram_ram_4(0), A2 => gl_ram_n_91, ZN => gl_ram_n_162);
  gl_ram_g56524 : ND2D2BWP7T port map(A1 => gl_ram_ram_87(1), A2 => gl_ram_n_92, ZN => gl_ram_n_161);
  gl_ram_g56526 : ND2D2BWP7T port map(A1 => gl_ram_ram_84(1), A2 => gl_ram_n_91, ZN => gl_ram_n_159);
  gl_ram_g56528 : ND2D2BWP7T port map(A1 => gl_ram_ram_83(1), A2 => gl_ram_n_87, ZN => gl_ram_n_157);
  gl_ram_g56529 : ND2D2BWP7T port map(A1 => gl_ram_ram_21(2), A2 => gl_ram_n_90, ZN => gl_ram_n_156);
  gl_ram_g56532 : ND2D2BWP7T port map(A1 => gl_ram_ram_95(1), A2 => gl_ram_n_92, ZN => gl_ram_n_153);
  gl_ram_g56535 : ND2D2BWP7T port map(A1 => gl_ram_ram_92(1), A2 => gl_ram_n_91, ZN => gl_ram_n_150);
  gl_ram_g56537 : ND2D2BWP7T port map(A1 => gl_ram_ram_90(1), A2 => gl_ram_n_86, ZN => gl_ram_n_148);
  gl_ram_g56539 : ND2D2BWP7T port map(A1 => gl_ram_ram_63(1), A2 => gl_ram_n_92, ZN => gl_ram_n_146);
  gl_ram_g56540 : CKND2D3BWP7T port map(A1 => gl_ram_ram_60(1), A2 => gl_ram_n_91, ZN => gl_ram_n_145);
  gl_ram_g56542 : ND2D2BWP7T port map(A1 => gl_ram_ram_62(1), A2 => gl_ram_n_93, ZN => gl_ram_n_143);
  gl_ram_g56548 : ND2D2BWP7T port map(A1 => gl_ram_ram_47(1), A2 => gl_ram_n_92, ZN => gl_ram_n_137);
  gl_ram_g56550 : ND2D2BWP7T port map(A1 => gl_ram_ram_44(1), A2 => gl_ram_n_91, ZN => gl_ram_n_135);
  gl_ram_g56553 : ND2D2BWP7T port map(A1 => gl_ram_ram_41(1), A2 => gl_ram_n_88, ZN => gl_ram_n_132);
  gl_ram_g56554 : ND2D1P5BWP7T port map(A1 => gl_ram_ram_43(1), A2 => gl_ram_n_87, ZN => gl_ram_n_131);
  gl_ram_g56557 : ND2D2BWP7T port map(A1 => gl_ram_ram_30(1), A2 => gl_ram_n_93, ZN => gl_ram_n_128);
  gl_ram_g56558 : ND2D2BWP7T port map(A1 => gl_ram_ram_31(1), A2 => gl_ram_n_92, ZN => gl_ram_n_127);
  gl_ram_g56559 : ND2D2BWP7T port map(A1 => gl_ram_ram_28(1), A2 => gl_ram_n_91, ZN => gl_ram_n_126);
  gl_ram_g56560 : CKND2D2BWP7T port map(A1 => gl_ram_ram_26(1), A2 => gl_ram_n_86, ZN => gl_ram_n_125);
  gl_ram_g56561 : ND2D2BWP7T port map(A1 => gl_ram_ram_25(1), A2 => gl_ram_n_88, ZN => gl_ram_n_124);
  gl_ram_g56563 : ND2D2BWP7T port map(A1 => gl_ram_ram_27(1), A2 => gl_ram_n_87, ZN => gl_ram_n_122);
  gl_ram_g56564 : ND2D2BWP7T port map(A1 => gl_ram_ram_39(1), A2 => gl_ram_n_92, ZN => gl_ram_n_121);
  gl_ram_g56565 : ND2D2BWP7T port map(A1 => gl_ram_ram_37(1), A2 => gl_ram_n_90, ZN => gl_ram_n_120);
  gl_ram_g56567 : ND2D2BWP7T port map(A1 => gl_ram_ram_36(1), A2 => gl_ram_n_91, ZN => gl_ram_n_118);
  gl_ram_g56569 : CKND2D2BWP7T port map(A1 => gl_ram_ram_34(1), A2 => gl_ram_n_86, ZN => gl_ram_n_116);
  gl_ram_g56572 : MAOI222D0BWP7T port map(A => gl_ram_y_grid(4), B => gl_ram_x_grid(4), C => gl_ram_y_grid(2), ZN => gl_ram_n_113);
  gl_ram_g56573 : ND2D2BWP7T port map(A1 => gl_ram_n_88, A2 => gl_ram_n_95, ZN => gl_ram_n_259);
  gl_ram_g56574 : ND2D2BWP7T port map(A1 => gl_ram_n_86, A2 => gl_ram_n_95, ZN => gl_ram_n_258);
  gl_ram_g56577 : AN2D2BWP7T port map(A1 => gl_ram_n_106, A2 => gl_ram_n_110, Z => gl_ram_n_256);
  gl_ram_g56581 : INVD5BWP7T port map(I => gl_ram_n_95, ZN => gl_ram_n_94);
  gl_ram_g56584 : OAI21D0BWP7T port map(A1 => gl_ram_n_1311, A2 => gl_ram_n_16, B => gl_ram_n_24, ZN => gl_ram_n_85);
  gl_ram_g56585 : ND2D1BWP7T port map(A1 => gl_ram_n_22, A2 => sig_output_color(0), ZN => gl_ram_n_112);
  gl_ram_g56586 : ND2D1BWP7T port map(A1 => gl_ram_n_22, A2 => sig_output_color(2), ZN => gl_ram_n_111);
  gl_ram_g56587 : ND2D1BWP7T port map(A1 => gl_ram_n_22, A2 => sig_output_color(1), ZN => gl_ram_n_110);
  gl_ram_g56588 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1244, A3 => FE_PHN347_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_780);
  gl_ram_g56589 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1246, A3 => FE_PHN289_gl_ram_n_1111, ZN => gl_ram_n_781);
  gl_ram_g56590 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1252, A3 => FE_PHN289_gl_ram_n_1111, ZN => gl_ram_n_784);
  gl_ram_g56591 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1254, A3 => FE_PHN289_gl_ram_n_1111, ZN => gl_ram_n_785);
  gl_ram_g56592 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1308, A3 => FE_PHN346_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_812);
  gl_ram_g56593 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1256, A3 => FE_PHN289_gl_ram_n_1111, ZN => gl_ram_n_786);
  gl_ram_g56594 : NR2D1P5BWP7T port map(A1 => gl_ram_n_22, A2 => gl_ram_ram_position(6), ZN => gl_ram_n_109);
  gl_ram_g56595 : IND2D4BWP7T port map(A1 => gl_ram_n_27, B1 => gl_ram_ram_position(4), ZN => gl_ram_n_108);
  gl_ram_g56596 : OR2D2BWP7T port map(A1 => gl_ram_n_27, A2 => gl_ram_ram_position(4), Z => gl_ram_n_107);
  gl_ram_g56598 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1248, A3 => FE_PHN289_gl_ram_n_1111, ZN => gl_ram_n_782);
  gl_ram_g56599 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1260, A3 => FE_PHN289_gl_ram_n_1111, ZN => gl_ram_n_788);
  gl_ram_g56600 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1250, A3 => FE_PHN289_gl_ram_n_1111, ZN => gl_ram_n_783);
  gl_ram_g56601 : ND2D1BWP7T port map(A1 => gl_ram_n_21, A2 => gl_ram_ram_position(6), ZN => gl_ram_n_106);
  gl_ram_g56602 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1268, A3 => FE_PHN325_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_792);
  gl_ram_g56603 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1258, A3 => FE_PHN289_gl_ram_n_1111, ZN => gl_ram_n_787);
  gl_ram_g56604 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1284, A3 => FE_PHN336_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_800);
  gl_ram_g56605 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1236, A3 => FE_PHN289_gl_ram_n_1111, ZN => gl_ram_n_776);
  gl_ram_g56606 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1270, A3 => FE_PHN344_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_793);
  gl_ram_g56607 : ND3D0BWP7T port map(A1 => CTS_345, A2 => gl_ram_n_1134, A3 => FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_105);
  gl_ram_g56608 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1304, A3 => FE_PHN339_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_810);
  gl_ram_g56609 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1302, A3 => FE_PHN348_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_809);
  gl_ram_g56610 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1298, A3 => FE_PHN339_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_807);
  gl_ram_g56611 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1296, A3 => FE_PHN339_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_806);
  gl_ram_g56612 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1294, A3 => FE_PHN339_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_805);
  gl_ram_g56613 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1292, A3 => FE_PHN336_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_804);
  gl_ram_g56614 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1290, A3 => FE_PHN336_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_803);
  gl_ram_g56615 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1288, A3 => FE_PHN345_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_802);
  gl_ram_g56616 : ND3D0BWP7T port map(A1 => CTS_344, A2 => gl_ram_n_1112, A3 => FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_103);
  gl_ram_g56617 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1286, A3 => FE_PHN336_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_801);
  gl_ram_g56618 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1282, A3 => FE_PHN336_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_799);
  gl_ram_g56619 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1280, A3 => FE_PHN336_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_798);
  gl_ram_g56620 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1278, A3 => FE_PHN336_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_797);
  gl_ram_g56621 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1234, A3 => FE_PHN289_gl_ram_n_1111, ZN => gl_ram_n_775);
  gl_ram_g56622 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1120, A3 => FE_PHN338_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_741);
  gl_ram_g56623 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1276, A3 => FE_PHN344_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_796);
  gl_ram_g56624 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1118, A3 => FE_PHN338_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_740);
  gl_ram_g56625 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1274, A3 => FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_795);
  gl_ram_g56626 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1272, A3 => FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_794);
  gl_ram_g56627 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1122, A3 => FE_PHN338_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_742);
  gl_ram_g56628 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1266, A3 => FE_PHN336_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_791);
  gl_ram_g56629 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1130, A3 => FE_PHN338_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_746);
  gl_ram_g56630 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1264, A3 => FE_PHN325_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_790);
  gl_ram_g56631 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1262, A3 => FE_PHN336_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_789);
  gl_ram_g56632 : ND3D0BWP7T port map(A1 => CTS_344, A2 => gl_ram_n_1156, A3 => FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_101);
  gl_ram_g56633 : ND2D6BWP7T port map(A1 => gl_ram_n_26, A2 => gl_ram_ram_position(4), ZN => gl_ram_n_99);
  gl_ram_g56634 : IND2D2BWP7T port map(A1 => gl_ram_ram_position(4), B1 => gl_ram_n_26, ZN => gl_ram_n_98);
  gl_ram_g56635 : ND2D6BWP7T port map(A1 => gl_ram_n_33, A2 => gl_ram_ram_position(4), ZN => gl_ram_n_97);
  gl_ram_g56636 : IND2D4BWP7T port map(A1 => gl_ram_ram_position(4), B1 => gl_ram_n_33, ZN => gl_ram_n_96);
  gl_ram_g56637 : NR2D0BWP7T port map(A1 => gl_ram_n_25, A2 => gl_ram_ram_position(4), ZN => gl_ram_n_95);
  gl_ram_g56638 : CKAN2D8BWP7T port map(A1 => gl_ram_n_32, A2 => gl_ram_ram_position(2), Z => gl_ram_n_93);
  gl_ram_g56639 : CKAN2D8BWP7T port map(A1 => gl_ram_n_29, A2 => gl_ram_ram_position(2), Z => gl_ram_n_92);
  gl_ram_g56640 : AN2D4BWP7T port map(A1 => gl_ram_n_31, A2 => gl_ram_ram_position(2), Z => gl_ram_n_91);
  gl_ram_g56641 : CKAN2D8BWP7T port map(A1 => gl_ram_n_30, A2 => gl_ram_ram_position(2), Z => gl_ram_n_90);
  gl_ram_g56642 : AN2D4BWP7T port map(A1 => gl_ram_n_31, A2 => gl_ram_n_17, Z => gl_ram_n_89);
  gl_ram_g56643 : AN2D4BWP7T port map(A1 => gl_ram_n_30, A2 => gl_ram_n_17, Z => gl_ram_n_88);
  gl_ram_g56644 : NR2D5BWP7T port map(A1 => gl_ram_n_28, A2 => gl_ram_ram_position(2), ZN => gl_ram_n_87);
  gl_ram_g56645 : AN2D4BWP7T port map(A1 => gl_ram_n_32, A2 => gl_ram_n_17, Z => gl_ram_n_86);
  gl_ram_g56670 : IOA21D0BWP7T port map(A1 => sig_logic_y(0), A2 => sig_logic_y(1), B => gl_ram_n_23, ZN => gl_ram_n_35);
  gl_ram_g56671 : MOAI22D0BWP7T port map(A1 => FE_PHN505_sig_logic_x_0, A2 => sig_logic_x(1), B1 => FE_PHN505_sig_logic_x_0, B2 => sig_logic_x(1), ZN => gl_ram_n_34);
  gl_ram_g56672 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1240, A3 => FE_PHN305_gl_ram_n_1111, ZN => gl_ram_n_778);
  gl_ram_g56673 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1238, A3 => FE_PHN340_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_777);
  gl_ram_g56674 : ND3D0BWP7T port map(A1 => CTS_344, A2 => gl_ram_n_1142, A3 => FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_84);
  gl_ram_g56675 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1232, A3 => FE_PHN289_gl_ram_n_1111, ZN => gl_ram_n_774);
  gl_ram_g56676 : ND3D0BWP7T port map(A1 => CTS_345, A2 => gl_ram_n_1146, A3 => FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_82);
  gl_ram_g56677 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1230, A3 => FE_PHN289_gl_ram_n_1111, ZN => gl_ram_n_773);
  gl_ram_g56678 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1228, A3 => FE_PHN337_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_772);
  gl_ram_g56679 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1226, A3 => FE_PHN309_gl_ram_n_1111, ZN => gl_ram_n_771);
  gl_ram_g56680 : ND3D0BWP7T port map(A1 => CTS_344, A2 => gl_ram_n_1150, A3 => FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_80);
  gl_ram_g56681 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1224, A3 => FE_PHN303_gl_ram_n_1111, ZN => gl_ram_n_770);
  gl_ram_g56682 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1222, A3 => FE_PHN337_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_769);
  gl_ram_g56683 : ND3D0BWP7T port map(A1 => CTS_345, A2 => gl_ram_n_1152, A3 => FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_78);
  gl_ram_g56684 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1218, A3 => FE_PHN300_gl_ram_n_1111, ZN => gl_ram_n_767);
  gl_ram_g56685 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1154, A3 => FE_PHN349_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_748);
  gl_ram_g56686 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1216, A3 => FE_PHN337_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_766);
  gl_ram_g56687 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1214, A3 => FE_PHN299_gl_ram_n_1111, ZN => gl_ram_n_765);
  gl_ram_g56688 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1212, A3 => FE_PHN341_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_764);
  gl_ram_g56689 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1210, A3 => FE_PHN341_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_763);
  gl_ram_g56690 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1300, A3 => FE_PHN339_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_808);
  gl_ram_g56691 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1208, A3 => FE_PHN341_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_762);
  gl_ram_g56692 : ND3D0BWP7T port map(A1 => CTS_344, A2 => gl_ram_n_1162, A3 => FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_76);
  gl_ram_g56693 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1202, A3 => FE_PHN341_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_759);
  gl_ram_g56694 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1200, A3 => FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_758);
  gl_ram_g56695 : ND3D0BWP7T port map(A1 => CTS_364, A2 => gl_ram_n_1166, A3 => FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_74);
  gl_ram_g56696 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1198, A3 => FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_757);
  gl_ram_g56697 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1196, A3 => FE_PHN289_gl_ram_n_1111, ZN => gl_ram_n_756);
  gl_ram_g56698 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1192, A3 => FE_PHN289_gl_ram_n_1111, ZN => gl_ram_n_754);
  gl_ram_g56699 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1190, A3 => FE_PHN289_gl_ram_n_1111, ZN => gl_ram_n_753);
  gl_ram_g56700 : ND3D0BWP7T port map(A1 => CTS_364, A2 => gl_ram_n_1172, A3 => FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_72);
  gl_ram_g56701 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1188, A3 => FE_PHN289_gl_ram_n_1111, ZN => gl_ram_n_752);
  gl_ram_g56702 : ND3D0BWP7T port map(A1 => CTS_345, A2 => gl_ram_n_1174, A3 => FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_70);
  gl_ram_g56703 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1184, A3 => FE_PHN289_gl_ram_n_1111, ZN => gl_ram_n_750);
  gl_ram_g56704 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1182, A3 => FE_PHN289_gl_ram_n_1111, ZN => gl_ram_n_749);
  gl_ram_g56705 : ND3D0BWP7T port map(A1 => CTS_345, A2 => gl_ram_n_1180, A3 => FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_68);
  gl_ram_g56706 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1186, A3 => FE_PHN289_gl_ram_n_1111, ZN => gl_ram_n_751);
  gl_ram_g56707 : ND3D0BWP7T port map(A1 => CTS_345, A2 => gl_ram_n_1176, A3 => FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_66);
  gl_ram_g56708 : ND3D0BWP7T port map(A1 => CTS_345, A2 => gl_ram_n_1178, A3 => FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_64);
  gl_ram_g56709 : ND3D0BWP7T port map(A1 => CTS_365, A2 => gl_ram_n_1168, A3 => FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_62);
  gl_ram_g56710 : ND3D0BWP7T port map(A1 => CTS_344, A2 => gl_ram_n_1164, A3 => FE_PHN335_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_60);
  gl_ram_g56711 : ND3D0BWP7T port map(A1 => CTS_345, A2 => gl_ram_n_1160, A3 => FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_58);
  gl_ram_g56712 : ND3D0BWP7T port map(A1 => CTS_345, A2 => gl_ram_n_1158, A3 => FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_56);
  gl_ram_g56713 : ND3D0BWP7T port map(A1 => CTS_364, A2 => gl_ram_n_1170, A3 => FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_54);
  gl_ram_g56714 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1194, A3 => FE_PHN289_gl_ram_n_1111, ZN => gl_ram_n_755);
  gl_ram_g56715 : ND3D0BWP7T port map(A1 => CTS_345, A2 => gl_ram_n_1148, A3 => FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_52);
  gl_ram_g56716 : ND3D0BWP7T port map(A1 => CTS_344, A2 => gl_ram_n_1144, A3 => FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_50);
  gl_ram_g56717 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1204, A3 => FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_760);
  gl_ram_g56718 : ND3D0BWP7T port map(A1 => CTS_344, A2 => gl_ram_n_1136, A3 => FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_48);
  gl_ram_g56719 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1206, A3 => FE_PHN341_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_761);
  gl_ram_g56720 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1132, A3 => FE_PHN342_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_747);
  gl_ram_g56721 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1128, A3 => FE_PHN338_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_745);
  gl_ram_g56722 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1126, A3 => FE_PHN342_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_744);
  gl_ram_g56723 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1124, A3 => FE_PHN338_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_743);
  gl_ram_g56724 : ND3D0BWP7T port map(A1 => CTS_364, A2 => gl_ram_n_1116, A3 => FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_46);
  gl_ram_g56725 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1220, A3 => FE_PHN317_gl_ram_n_1111, ZN => gl_ram_n_768);
  gl_ram_g56726 : ND3D0BWP7T port map(A1 => CTS_364, A2 => gl_ram_n_1110, A3 => FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_44);
  gl_ram_g56727 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1242, A3 => FE_PHN343_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_779);
  gl_ram_g56728 : ND3D0BWP7T port map(A1 => CTS_289, A2 => gl_ram_n_1306, A3 => FE_PHN339_FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_811);
  gl_ram_g56729 : ND3D0BWP7T port map(A1 => CTS_344, A2 => gl_ram_n_1114, A3 => FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_42);
  gl_ram_g56730 : ND3D0BWP7T port map(A1 => CTS_364, A2 => gl_ram_n_1140, A3 => FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_40);
  gl_ram_g56731 : ND3D0BWP7T port map(A1 => CTS_344, A2 => gl_ram_n_1138, A3 => FE_OFN4_gl_ram_n_1111, ZN => gl_ram_n_38);
  gl_ram_g56732 : XNR2D1BWP7T port map(A1 => gl_ram_x_grid(4), A2 => gl_ram_y_grid(4), ZN => gl_ram_n_36);
  gl_ram_g56734 : INR2D0BWP7T port map(A1 => gl_ram_ram_position(3), B1 => gl_ram_ram_position(5), ZN => gl_ram_n_33);
  gl_ram_g56735 : INR2D0BWP7T port map(A1 => gl_ram_ram_position(1), B1 => gl_ram_ram_position(0), ZN => gl_ram_n_32);
  gl_ram_g56736 : NR2D0BWP7T port map(A1 => gl_ram_ram_position(1), A2 => gl_ram_ram_position(0), ZN => gl_ram_n_31);
  gl_ram_g56740 : CKND1BWP7T port map(I => gl_ram_n_28, ZN => gl_ram_n_29);
  gl_ram_g56742 : INVD1BWP7T port map(I => gl_ram_n_21, ZN => gl_ram_n_22);
  gl_ram_g56743 : INR2D0BWP7T port map(A1 => gl_ram_ram_position(0), B1 => gl_ram_ram_position(1), ZN => gl_ram_n_30);
  gl_ram_g56744 : ND2D0BWP7T port map(A1 => gl_ram_ram_position(1), A2 => gl_ram_ram_position(0), ZN => gl_ram_n_28);
  gl_ram_g56745 : ND2D0BWP7T port map(A1 => gl_ram_ram_position(5), A2 => gl_ram_ram_position(3), ZN => gl_ram_n_27);
  gl_ram_g56746 : NR2D0BWP7T port map(A1 => gl_ram_ram_position(5), A2 => gl_ram_ram_position(3), ZN => gl_ram_n_26);
  gl_ram_g56747 : IND2D0BWP7T port map(A1 => gl_ram_ram_position(3), B1 => gl_ram_ram_position(5), ZN => gl_ram_n_25);
  gl_ram_g56748 : ND2D0BWP7T port map(A1 => gl_ram_n_1311, A2 => gl_ram_n_16, ZN => gl_ram_n_24);
  gl_ram_g56749 : IND2D0BWP7T port map(A1 => sig_logic_y(1), B1 => gl_ram_n_19, ZN => gl_ram_n_23);
  gl_ram_g56750 : ND2D1BWP7T port map(A1 => sig_rescount, A2 => sig_draw, ZN => gl_ram_n_21);
  gl_ram_g56766 : CKND1BWP7T port map(I => sig_logic_y(0), ZN => gl_ram_n_19);
  gl_ram_g56767 : CKND1BWP7T port map(I => FE_PHN505_sig_logic_x_0, ZN => gl_ram_n_18);
  gl_ram_g56768 : INVD0BWP7T port map(I => gl_ram_ram_position(2), ZN => gl_ram_n_17);
  gl_ram_g56769 : CKND1BWP7T port map(I => FE_PHN315_sig_logic_x_2, ZN => gl_ram_n_16);
  gl_ram_g56782 : INR2D1BWP7T port map(A1 => gl_ram_n_89, B1 => gl_ram_n_94, ZN => gl_ram_n_6);
  gl_ram_g56783 : INR2D1BWP7T port map(A1 => gl_ram_n_87, B1 => gl_ram_n_94, ZN => gl_ram_n_5);
  gl_ram_g56784 : IND2D2BWP7T port map(A1 => gl_ram_n_25, B1 => gl_ram_ram_position(4), ZN => gl_ram_n_4);
  gl_ram_g56786 : INR2D4BWP7T port map(A1 => gl_ram_ram_98(1), B1 => gl_ram_n_258, ZN => gl_ram_n_2);
  gl_ram_ram_reg_28_1 : LND1BWP7T port map(D => gl_ram_n_1446, EN => gl_ram_n_784, Q => gl_ram_ram_28(1), QN => UNCONNECTED);
  gl_ram_ram_reg_28_2 : LND2BWP7T port map(D => FE_OCPN3_gl_ram_n_1448, EN => gl_ram_n_784, Q => gl_ram_ram_28(2), QN => UNCONNECTED0);
  gl_ram_g56805 : ND2D6BWP7T port map(A1 => gl_ram_n_727, A2 => gl_ram_n_732, ZN => gl_ram_n_1436);
  gl_ram_g55934_dup : ND2D5BWP7T port map(A1 => gl_ram_n_732, A2 => gl_ram_n_727, ZN => gl_ram_n_1437);
  gl_ram_ram_reg_57_0 : LND1BWP7T port map(D => gl_ram_n_1437, EN => gl_ram_n_755, Q => gl_ram_ram_57(0), QN => UNCONNECTED1);
  gl_ram_ram_reg_58_0 : LND1BWP7T port map(D => gl_ram_n_1436, EN => gl_ram_n_754, Q => gl_ram_ram_58(0), QN => UNCONNECTED2);
  gl_ram_ram_reg_25_0 : LND1BWP7T port map(D => gl_ram_n_1436, EN => gl_ram_n_787, Q => gl_ram_ram_25(0), QN => UNCONNECTED3);
  gl_ram_g56829 : NR2XD2BWP7T port map(A1 => gl_ram_n_1438, A2 => gl_ram_n_475, ZN => gl_ram_n_1439);
  gl_ram_ram_reg_63_0 : LND2BWP7T port map(D => gl_ram_n_1437, EN => gl_ram_n_749, Q => gl_ram_ram_63(0), QN => UNCONNECTED4);
  gl_ram_ram_reg_26_0 : LND1BWP7T port map(D => gl_ram_n_1436, EN => gl_ram_n_786, Q => gl_ram_ram_26(0), QN => UNCONNECTED5);
  gl_ram_ram_reg_61_0 : LND1BWP7T port map(D => gl_ram_n_1436, EN => gl_ram_n_751, Q => gl_ram_ram_61(0), QN => UNCONNECTED6);
  gl_ram_ram_reg_9_0 : LND1BWP7T port map(D => gl_ram_n_736, EN => gl_ram_n_803, Q => gl_ram_ram_9(0), QN => UNCONNECTED7);
  gl_ram_ram_reg_57_1 : LND1BWP7T port map(D => gl_ram_n_735, EN => gl_ram_n_755, Q => gl_ram_ram_57(1), QN => UNCONNECTED8);
  gl_ram_ram_reg_57_2 : LND2BWP7T port map(D => gl_ram_n_739, EN => gl_ram_n_755, Q => gl_ram_ram_57(2), QN => UNCONNECTED9);
  gl_ram_fopt : INVD4BWP7T port map(I => gl_ram_ram_97(0), ZN => gl_ram_n_1440);
  gl_ram_ram_reg_17_0 : LND1BWP7T port map(D => gl_ram_n_736, EN => gl_ram_n_795, Q => gl_ram_ram_17(0), QN => UNCONNECTED10);
  gl_ram_ram_reg_58_1 : LND1BWP7T port map(D => gl_ram_n_735, EN => gl_ram_n_754, Q => gl_ram_ram_58(1), QN => UNCONNECTED11);
  gl_ram_ram_reg_58_2 : LND1BWP7T port map(D => gl_ram_n_739, EN => gl_ram_n_754, Q => gl_ram_ram_58(2), QN => UNCONNECTED12);
  gl_ram_ram_reg_28_0 : LND1BWP7T port map(D => gl_ram_n_1437, EN => gl_ram_n_784, Q => gl_ram_ram_28(0), QN => UNCONNECTED13);
  gl_ram_ram_reg_30_0 : LND1BWP7T port map(D => gl_ram_n_1437, EN => gl_ram_n_782, Q => gl_ram_ram_30(0), QN => UNCONNECTED14);
  gl_ram_g56869 : NR2XD2BWP7T port map(A1 => gl_ram_n_1444, A2 => gl_ram_n_1521, ZN => gl_ram_n_1445);
  gl_ram_g56870 : IOA21D2BWP7T port map(A1 => gl_ram_ram_16(0), A2 => gl_ram_n_89, B => gl_ram_n_178, ZN => gl_ram_n_1444);
  gl_ram_g56871 : ND2D5BWP7T port map(A1 => gl_ram_n_731, A2 => gl_ram_n_726, ZN => gl_ram_n_1446);
  gl_ram_g55937_dup : ND2D5BWP7T port map(A1 => gl_ram_n_731, A2 => gl_ram_n_726, ZN => gl_ram_n_1447);
  gl_ram_g56872 : ND2D4BWP7T port map(A1 => gl_ram_n_733, A2 => gl_ram_n_728, ZN => gl_ram_n_1448);
  gl_ram_g56904 : AN2D4BWP7T port map(A1 => gl_ram_ram_99(1), A2 => gl_ram_n_5, Z => gl_ram_n_1450);
  gl_ram_g56905 : AOI22D2BWP7T port map(A1 => gl_ram_ram_96(0), A2 => gl_ram_n_6, B1 => gl_ram_ram_99(0), B2 => gl_ram_n_5, ZN => gl_ram_n_1451);
  gl_ram_g56909 : IOA21D2BWP7T port map(A1 => gl_ram_ram_22(1), A2 => gl_ram_n_93, B => gl_ram_n_391, ZN => gl_ram_n_1455);
  gl_ram_g56910 : IOA21D2BWP7T port map(A1 => gl_ram_ram_16(1), A2 => gl_ram_n_89, B => gl_ram_n_388, ZN => gl_ram_n_1456);
  gl_ram_g56911 : IOA21D2BWP7T port map(A1 => gl_ram_ram_54(1), A2 => gl_ram_n_93, B => gl_ram_n_381, ZN => gl_ram_n_1457);
  gl_ram_g56912 : IOA21D2BWP7T port map(A1 => gl_ram_ram_48(1), A2 => gl_ram_n_89, B => gl_ram_n_378, ZN => gl_ram_n_1458);
  gl_ram_g56914 : IOA21D2BWP7T port map(A1 => gl_ram_ram_6(1), A2 => gl_ram_n_93, B => gl_ram_n_373, ZN => gl_ram_n_1460);
  gl_ram_g56915 : IOA21D2BWP7T port map(A1 => gl_ram_ram_1(1), A2 => gl_ram_n_88, B => gl_ram_n_371, ZN => gl_ram_n_1461);
  gl_ram_g56916 : IOA21D2BWP7T port map(A1 => gl_ram_ram_0(1), A2 => gl_ram_n_89, B => gl_ram_n_387, ZN => gl_ram_n_1462);
  gl_ram_g56920 : IOA21D2BWP7T port map(A1 => gl_ram_ram_72(2), A2 => gl_ram_n_89, B => gl_ram_n_361, ZN => gl_ram_n_1466);
  gl_ram_g56922 : IOA21D2BWP7T port map(A1 => gl_ram_ram_65(2), A2 => gl_ram_n_88, B => gl_ram_n_354, ZN => gl_ram_n_1468);
  gl_ram_g56923 : IOA21D2BWP7T port map(A1 => gl_ram_ram_64(2), A2 => gl_ram_n_89, B => gl_ram_n_353, ZN => gl_ram_n_1469);
  gl_ram_g56926 : IOA21D2BWP7T port map(A1 => gl_ram_ram_81(2), A2 => gl_ram_n_88, B => gl_ram_n_345, ZN => gl_ram_n_1472);
  gl_ram_g56927 : IOA21D2BWP7T port map(A1 => gl_ram_ram_93(2), A2 => gl_ram_n_90, B => gl_ram_n_343, ZN => gl_ram_n_1473);
  gl_ram_g56935 : IOA21D2BWP7T port map(A1 => gl_ram_ram_42(2), A2 => gl_ram_n_86, B => gl_ram_n_322, ZN => gl_ram_n_1481);
  gl_ram_g56938 : IOA21D2BWP7T port map(A1 => gl_ram_ram_25(2), A2 => gl_ram_n_88, B => gl_ram_n_315, ZN => gl_ram_n_1484);
  gl_ram_g56939 : IOA21D2BWP7T port map(A1 => gl_ram_ram_38(2), A2 => gl_ram_n_93, B => gl_ram_n_360, ZN => gl_ram_n_1485);
  gl_ram_g56940 : IOA21D2BWP7T port map(A1 => gl_ram_ram_33(2), A2 => gl_ram_n_88, B => gl_ram_n_307, ZN => gl_ram_n_1486);
  gl_ram_g56942 : IOA21D2BWP7T port map(A1 => gl_ram_ram_13(2), A2 => gl_ram_n_90, B => gl_ram_n_303, ZN => gl_ram_n_1488);
  gl_ram_g56943 : IOA21D2BWP7T port map(A1 => gl_ram_ram_9(2), A2 => gl_ram_n_88, B => gl_ram_n_299, ZN => gl_ram_n_1489);
  gl_ram_g56944 : IOA21D2BWP7T port map(A1 => gl_ram_ram_22(2), A2 => gl_ram_n_93, B => gl_ram_n_292, ZN => gl_ram_n_1490);
  gl_ram_g56945 : IOA21D2BWP7T port map(A1 => gl_ram_ram_13(0), A2 => gl_ram_n_90, B => gl_ram_n_188, ZN => gl_ram_n_1491);
  gl_ram_g56946 : IOA21D2BWP7T port map(A1 => gl_ram_ram_48(2), A2 => gl_ram_n_89, B => gl_ram_n_279, ZN => gl_ram_n_1492);
  gl_ram_g56947 : IOA21D2BWP7T port map(A1 => gl_ram_ram_5(2), A2 => gl_ram_n_90, B => gl_ram_n_276, ZN => gl_ram_n_1493);
  gl_ram_g56948 : IOA21D2BWP7T port map(A1 => gl_ram_ram_72(0), A2 => gl_ram_n_89, B => gl_ram_n_277, ZN => gl_ram_n_1494);
  gl_ram_g56950 : IOA21D2BWP7T port map(A1 => gl_ram_ram_0(2), A2 => gl_ram_n_89, B => gl_ram_n_271, ZN => gl_ram_n_1496);
  gl_ram_g56951 : IOA21D2BWP7T port map(A1 => gl_ram_ram_1(2), A2 => gl_ram_n_88, B => gl_ram_n_273, ZN => gl_ram_n_1497);
  gl_ram_g56954 : IOA21D2BWP7T port map(A1 => gl_ram_ram_69(1), A2 => gl_ram_n_90, B => gl_ram_n_267, ZN => gl_ram_n_1500);
  gl_ram_g56955 : IOA21D2BWP7T port map(A1 => gl_ram_ram_80(0), A2 => gl_ram_n_89, B => gl_ram_n_249, ZN => gl_ram_n_1501);
  gl_ram_g56956 : IOA21D2BWP7T port map(A1 => gl_ram_ram_77(1), A2 => gl_ram_n_90, B => gl_ram_n_243, ZN => gl_ram_n_1502);
  gl_ram_g56957 : IOA21D2BWP7T port map(A1 => gl_ram_ram_89(0), A2 => gl_ram_n_88, B => gl_ram_n_232, ZN => gl_ram_n_1503);
  gl_ram_g56961 : IOA21D2BWP7T port map(A1 => gl_ram_ram_62(0), A2 => gl_ram_n_93, B => gl_ram_n_229, ZN => gl_ram_n_1507);
  gl_ram_g56962 : IOA21D2BWP7T port map(A1 => gl_ram_ram_45(0), A2 => gl_ram_n_90, B => gl_ram_n_220, ZN => gl_ram_n_1508);
  gl_ram_g56965 : IOA21D2BWP7T port map(A1 => gl_ram_ram_29(0), A2 => gl_ram_n_90, B => gl_ram_n_205, ZN => gl_ram_n_1511);
  gl_ram_g56968 : IOA21D2BWP7T port map(A1 => gl_ram_ram_38(0), A2 => gl_ram_n_93, B => gl_ram_n_174, ZN => gl_ram_n_1514);
  gl_ram_g56971 : IOA21D2BWP7T port map(A1 => gl_ram_ram_54(2), A2 => gl_ram_n_93, B => gl_ram_n_283, ZN => gl_ram_n_1517);
  gl_ram_g56972 : IOA21D2BWP7T port map(A1 => gl_ram_ram_9(0), A2 => gl_ram_n_88, B => gl_ram_n_185, ZN => gl_ram_n_1518);
  gl_ram_g56973 : IOA21D2BWP7T port map(A1 => gl_ram_ram_8(0), A2 => gl_ram_n_89, B => gl_ram_n_183, ZN => gl_ram_n_1519);
  gl_ram_g56974 : IOA21D2BWP7T port map(A1 => gl_ram_ram_22(0), A2 => gl_ram_n_93, B => gl_ram_n_179, ZN => gl_ram_n_1520);
  gl_ram_g56975 : IOA21D2BWP7T port map(A1 => gl_ram_ram_17(0), A2 => gl_ram_n_88, B => gl_ram_n_192, ZN => gl_ram_n_1521);
  gl_ram_g56980 : IOA21D2BWP7T port map(A1 => gl_ram_ram_78(1), A2 => gl_ram_n_93, B => gl_ram_n_269, ZN => gl_ram_n_1526);
  gl_ram_g56981 : IOA21D2BWP7T port map(A1 => gl_ram_ram_72(1), A2 => gl_ram_n_89, B => gl_ram_n_168, ZN => gl_ram_n_1527);
  gl_ram_g56982 : IOA21D2BWP7T port map(A1 => gl_ram_ram_64(1), A2 => gl_ram_n_89, B => gl_ram_n_166, ZN => gl_ram_n_1528);
  gl_ram_g56983 : IOA21D2BWP7T port map(A1 => gl_ram_ram_70(1), A2 => gl_ram_n_93, B => gl_ram_n_163, ZN => gl_ram_n_1529);
  gl_ram_g56984 : IOA21D2BWP7T port map(A1 => gl_ram_ram_65(1), A2 => gl_ram_n_88, B => gl_ram_n_245, ZN => gl_ram_n_1530);
  gl_ram_g56985 : IOA21D2BWP7T port map(A1 => gl_ram_ram_85(1), A2 => gl_ram_n_90, B => gl_ram_n_161, ZN => gl_ram_n_1531);
  gl_ram_g56986 : IOA21D2BWP7T port map(A1 => gl_ram_ram_80(1), A2 => gl_ram_n_89, B => gl_ram_n_157, ZN => gl_ram_n_1532);
  gl_ram_g56987 : IOA21D2BWP7T port map(A1 => gl_ram_ram_86(1), A2 => gl_ram_n_93, B => gl_ram_n_159, ZN => gl_ram_n_1533);
  gl_ram_g56988 : IOA21D2BWP7T port map(A1 => gl_ram_ram_93(1), A2 => gl_ram_n_90, B => gl_ram_n_153, ZN => gl_ram_n_1534);
  gl_ram_g56989 : IOA21D2BWP7T port map(A1 => gl_ram_ram_94(1), A2 => gl_ram_n_93, B => gl_ram_n_150, ZN => gl_ram_n_1535);
  gl_ram_g56990 : IOA21D2BWP7T port map(A1 => gl_ram_ram_89(1), A2 => gl_ram_n_88, B => gl_ram_n_148, ZN => gl_ram_n_1536);
  gl_ram_g56991 : IOA21D2BWP7T port map(A1 => gl_ram_ram_88(1), A2 => gl_ram_n_89, B => gl_ram_n_181, ZN => gl_ram_n_1537);
  gl_ram_g56994 : IOA21D2BWP7T port map(A1 => gl_ram_ram_45(1), A2 => gl_ram_n_90, B => gl_ram_n_137, ZN => gl_ram_n_1540);
  gl_ram_g56996 : IOA21D2BWP7T port map(A1 => gl_ram_ram_42(1), A2 => gl_ram_n_86, B => gl_ram_n_132, ZN => gl_ram_n_1542);
  gl_ram_g56997 : IOA21D2BWP7T port map(A1 => gl_ram_ram_40(1), A2 => gl_ram_n_89, B => gl_ram_n_131, ZN => gl_ram_n_1543);
  gl_ram_g56998 : IOA21D2BWP7T port map(A1 => gl_ram_ram_29(1), A2 => gl_ram_n_90, B => gl_ram_n_127, ZN => gl_ram_n_1544);
  gl_ram_g56999 : IOA21D2BWP7T port map(A1 => gl_ram_ram_24(1), A2 => gl_ram_n_89, B => gl_ram_n_122, ZN => gl_ram_n_1545);
  gl_ram_g57000 : IOA21D2BWP7T port map(A1 => gl_ram_ram_38(1), A2 => gl_ram_n_93, B => gl_ram_n_118, ZN => gl_ram_n_1546);
  gl_ram_g57001 : IOA21D2BWP7T port map(A1 => gl_ram_ram_32(1), A2 => gl_ram_n_89, B => gl_ram_n_240, ZN => gl_ram_n_1547);
  gl_ram_g57002 : IOA21D2BWP7T port map(A1 => gl_ram_ram_33(1), A2 => gl_ram_n_88, B => gl_ram_n_116, ZN => gl_ram_n_1548);
  gl_ram_ram_reg_12_0 : LND1BWP7T port map(D => gl_ram_n_736, EN => gl_ram_n_800, Q => gl_ram_ram_12(0), QN => UNCONNECTED15);
  gl_ram_g57007 : IOA21D2BWP7T port map(A1 => gl_ram_ram_69(2), A2 => gl_ram_n_90, B => gl_ram_n_359, ZN => gl_ram_n_1551);
  gl_ram_g57008 : IOA21D2BWP7T port map(A1 => gl_ram_ram_64(0), A2 => gl_ram_n_89, B => gl_ram_n_304, ZN => gl_ram_n_1552);
  gl_ram_ram_reg_33_0 : LNQD1BWP7T port map(D => gl_ram_n_1437, EN => gl_ram_n_779, Q => gl_ram_ram_33(0));
  gl_ram_ram_reg_41_0 : LNQD2BWP7T port map(D => gl_ram_n_1437, EN => gl_ram_n_771, Q => gl_ram_ram_41(0));
  gl_ram_ram_reg_41_1 : LNQD1BWP7T port map(D => gl_ram_n_1447, EN => gl_ram_n_771, Q => gl_ram_ram_41(1));
  gl_ram_ram_reg_30_1 : LNQD1BWP7T port map(D => gl_ram_n_1447, EN => gl_ram_n_782, Q => gl_ram_ram_30(1));
  gl_ram_ram_reg_31_1 : LNQD1BWP7T port map(D => gl_ram_n_1446, EN => gl_ram_n_781, Q => gl_ram_ram_31(1));
  gl_ram_ram_reg_41_2 : LNQD1BWP7T port map(D => gl_ram_n_1449, EN => gl_ram_n_771, Q => gl_ram_ram_41(2));
  gl_ram_ram_reg_30_2 : LNQD2BWP7T port map(D => FE_OCPN3_gl_ram_n_1448, EN => gl_ram_n_782, Q => gl_ram_ram_30(2));
  gl_ram_ram_reg_31_2 : LNQD2BWP7T port map(D => FE_OCPN3_gl_ram_n_1448, EN => gl_ram_n_781, Q => gl_ram_ram_31(2));
  ml_ms_g754 : OR2D1BWP7T port map(A1 => ml_ms_n_62, A2 => ml_ms_n_63, Z => FE_OFN33_clk15k_switch);
  ml_ms_g755 : INR2XD0BWP7T port map(A1 => ml_ms_sfsm_n_383, B1 => ml_ms_muxFSM, ZN => ml_ms_n_63);
  ml_ms_g757 : NR2XD0BWP7T port map(A1 => ml_ms_n_61, A2 => FE_PHN416_ml_ms_sfsm_state_0, ZN => ml_ms_n_62);
  ml_ms_g758 : CKAN2D1BWP7T port map(A1 => ml_ms_sfsm_state(1), A2 => FE_PHN416_ml_ms_sfsm_state_0, Z => ml_ms_sfsm_n_383);
  ml_ms_g760 : IND2D1BWP7T port map(A1 => ml_ms_sfsm_state(1), B1 => ml_ms_muxFSM, ZN => ml_ms_n_61);
  ml_ms_g2 : INR2D1BWP7T port map(A1 => ml_ms_n_61, B1 => FE_PHN416_ml_ms_sfsm_state_0, ZN => ml_ms_cntReset25M_send);
  ml_ms_sfsm_state_reg_0 : DFQD1BWP7T port map(CP => CTS_322, D => FE_PHN480_ml_ms_n_58, Q => ml_ms_sfsm_state(0));
  ml_ms_sr_new_new_data_reg_0 : DFQD1BWP7T port map(CP => CTS_288, D => FE_PHN460_ml_ms_n_30, Q => ml_ms_sr_new_new_data(0));
  ml_ms_sr_new_new_data_reg_1 : DFQD1BWP7T port map(CP => CTS_288, D => ml_ms_n_20, Q => ml_ms_sr_new_new_data(1));
  ml_ms_sr_new_new_data_reg_2 : DFQD1BWP7T port map(CP => CTS_288, D => ml_ms_n_19, Q => ml_ms_sr_new_new_data(2));
  ml_ms_sr_new_new_data_reg_3 : DFQD1BWP7T port map(CP => CTS_288, D => ml_ms_n_26, Q => ml_ms_sr_new_new_data(3));
  ml_ms_sr_new_new_data_reg_4 : DFQD1BWP7T port map(CP => CTS_288, D => ml_ms_n_25, Q => ml_ms_sr_new_new_data(4));
  ml_ms_sr_new_new_data_reg_5 : DFQD1BWP7T port map(CP => CTS_288, D => ml_ms_n_34, Q => ml_ms_sr_new_new_data(5));
  ml_ms_sr_new_new_data_reg_6 : DFQD1BWP7T port map(CP => CTS_288, D => FE_PHN462_ml_ms_n_24, Q => ml_ms_sr_new_new_data(6));
  ml_ms_sr_new_new_data_reg_7 : DFQD1BWP7T port map(CP => CTS_288, D => FE_PHN458_ml_ms_n_32, Q => ml_ms_sr_new_new_data(7));
  ml_ms_sr_new_new_data_reg_8 : DFQD1BWP7T port map(CP => CTS_288, D => FE_PHN463_ml_ms_n_31, Q => ml_ms_muxReg);
  ml_ms_g1847 : MOAI22D0BWP7T port map(A1 => ml_ms_n_45, A2 => ml_ms_n_10, B1 => ml_ms_n_59, B2 => FE_PHN425_ml_ms_mux_select, ZN => ml_ms_n_60);
  ml_ms_g1850 : OAI211D1BWP7T port map(A1 => ml_ms_n_8, A2 => ml_ms_n_47, B => ml_ms_n_55, C => ml_ms_n_52, ZN => ml_ms_n_59);
  ml_ms_g1851 : OAI211D1BWP7T port map(A1 => ml_ms_n_49, A2 => ml_ms_n_53, B => ml_ms_n_56, C => ml_ms_n_52, ZN => ml_ms_n_58);
  ml_ms_g1852 : OAI221D0BWP7T port map(A1 => ml_ms_n_53, A2 => ml_ms_n_50, B1 => ml_ms_n_0, B2 => ml_ms_n_8, C => ml_ms_n_51, ZN => ml_ms_n_57);
  ml_ms_g1854 : OAI21D0BWP7T port map(A1 => ml_ms_n_47, A2 => ml_ms_n_14, B => ml_ms_n_7, ZN => ml_ms_n_56);
  ml_ms_g1855 : IND3D1BWP7T port map(A1 => ml_ms_n_10, B1 => ml_ms_muxFSM, B2 => ml_ms_n_50, ZN => ml_ms_n_55);
  ml_ms_g1856 : MOAI22D0BWP7T port map(A1 => ml_ms_n_48, A2 => ml_ms_n_16, B1 => ml_ms_n_46, B2 => ml_ms_muxFSM, ZN => ml_ms_n_54);
  ml_ms_g1857 : IND3D1BWP7T port map(A1 => ml_ms_n_10, B1 => ml_ms_muxFSM, B2 => ml_ms_n_45, ZN => ml_ms_n_53);
  ml_ms_g1858 : IND3D1BWP7T port map(A1 => ml_ms_n_40, B1 => ml_ms_n_45, B2 => ml_ms_n_48, ZN => ml_ms_n_51);
  ml_ms_g1859 : IND3D1BWP7T port map(A1 => ml_ms_n_16, B1 => ml_ms_n_37, B2 => ml_ms_n_48, ZN => ml_ms_n_52);
  ml_ms_g1860 : INVD0BWP7T port map(I => ml_ms_n_50, ZN => ml_ms_n_49);
  ml_ms_g1861 : IAO21D0BWP7T port map(A1 => ml_ms_n_43, A2 => ml_ms_n_11, B => ml_ms_count25M(12), ZN => ml_ms_n_50);
  ml_ms_g1862 : IOA21D1BWP7T port map(A1 => ml_ms_n_42, A2 => ml_ms_n_18, B => ml_ms_sfsm_state(1), ZN => ml_ms_n_48);
  ml_ms_g1863 : AOI21D0BWP7T port map(A1 => ml_ms_n_44, A2 => FE_PHN416_ml_ms_sfsm_state_0, B => ml_ms_reset_send, ZN => ml_ms_n_46);
  ml_ms_g1864 : AOI211XD0BWP7T port map(A1 => ml_ms_sfsm_state(1), A2 => FE_PHN438_clk15k_in, B => ml_ms_n_41, C => ml_ms_n_1, ZN => ml_ms_n_47);
  ml_ms_g1865 : ND2D1BWP7T port map(A1 => ml_ms_n_44, A2 => ml_ms_muxFSM, ZN => ml_ms_n_45);
  ml_ms_g1866 : NR2XD0BWP7T port map(A1 => ml_ms_n_38, A2 => ml_ms_count25M(9), ZN => ml_ms_n_43);
  ml_ms_g1867 : OA31D1BWP7T port map(A1 => ml_ms_count25M(11), A2 => ml_ms_count25M(10), A3 => ml_ms_n_33, B => ml_ms_sfsm_state(1), Z => ml_ms_n_44);
  ml_ms_g1868 : OAI211D1BWP7T port map(A1 => ml_ms_n_17, A2 => ml_ms_n_36, B => ml_ms_count25M(11), C => ml_ms_count25M(9), ZN => ml_ms_n_42);
  ml_ms_g1869 : NR2D1BWP7T port map(A1 => ml_ms_n_39, A2 => ml_ms_sfsm_state(1), ZN => ml_ms_n_41);
  ml_ms_g1870 : OA22D0BWP7T port map(A1 => ml_ms_n_16, A2 => ml_ms_n_37, B1 => ml_ms_n_0, B2 => ml_ms_n_10, Z => ml_ms_n_40);
  ml_ms_g1871 : AOI21D0BWP7T port map(A1 => ml_ms_n_35, A2 => ml_ms_n_15, B => ml_ms_n_18, ZN => ml_ms_n_39);
  ml_ms_g1872 : AO211D0BWP7T port map(A1 => ml_ms_n_27, A2 => ml_ms_count25M(8), B => ml_ms_n_29, C => ml_ms_n_17, Z => ml_ms_n_38);
  ml_ms_g1877 : ND4D0BWP7T port map(A1 => ml_ms_n_12, A2 => ml_ms_count25M(8), A3 => ml_ms_count25M(9), A4 => ml_ms_count25M(12), ZN => ml_ms_n_37);
  ml_ms_g1878 : AN2D0BWP7T port map(A1 => ml_ms_n_29, A2 => ml_ms_count25M(3), Z => ml_ms_n_36);
  ml_ms_g1884 : OAI211D1BWP7T port map(A1 => ml_ms_count25M(3), A2 => ml_ms_n_3, B => ml_ms_n_5, C => ml_ms_count25M(5), ZN => ml_ms_n_35);
  ml_ms_g1885 : ND2D1BWP7T port map(A1 => ml_ms_n_28, A2 => ml_ms_n_22, ZN => FE_PHN464_ml_ms_n_34);
  ml_ms_g1886 : OAI21D0BWP7T port map(A1 => ml_ms_n_13, A2 => ml_ms_n_6, B => ml_ms_n_15, ZN => ml_ms_n_33);
  ml_ms_g1887 : ND2D1BWP7T port map(A1 => ml_ms_n_28, A2 => ml_ms_n_23, ZN => ml_ms_n_32);
  ml_ms_g1888 : ND2D1BWP7T port map(A1 => ml_ms_n_28, A2 => ml_ms_n_21, ZN => ml_ms_n_31);
  ml_ms_g1889 : IOA21D1BWP7T port map(A1 => ml_ms_n_4, A2 => ml_ms_sr_new_new_data(0), B => ml_ms_n_28, ZN => ml_ms_n_30);
  ml_ms_g1890 : AN4D0BWP7T port map(A1 => ml_ms_count25M(3), A2 => ml_ms_count25M(2), A3 => ml_ms_count25M(7), A4 => ml_ms_count25M(5), Z => ml_ms_n_27);
  ml_ms_g1891 : AO22D0BWP7T port map(A1 => ml_ms_n_4, A2 => ml_ms_sr_new_new_data(3), B1 => ml_ms_sr_new_new_data(2), B2 => ml_ms_n_9, Z => FE_PHN461_ml_ms_n_26);
  ml_ms_g1892 : AO22D0BWP7T port map(A1 => ml_ms_n_4, A2 => ml_ms_sr_new_new_data(4), B1 => ml_ms_sr_new_new_data(3), B2 => ml_ms_n_9, Z => FE_PHN465_ml_ms_n_25);
  ml_ms_g1893 : AN4D0BWP7T port map(A1 => FE_PHN437_ml_ms_count25M_4, A2 => ml_ms_count25M(8), A3 => ml_ms_count25M(7), A4 => ml_ms_count25M(5), Z => ml_ms_n_29);
  ml_ms_g1894 : OAI211D1BWP7T port map(A1 => ml_ms_muxFSM, A2 => ml_ms_sfsm_n_383, B => ml_ms_actBit, C => ml_ms_n_2, ZN => ml_ms_n_28);
  ml_ms_g1895 : AO22D0BWP7T port map(A1 => ml_ms_n_4, A2 => ml_ms_sr_new_new_data(6), B1 => ml_ms_sr_new_new_data(5), B2 => ml_ms_n_9, Z => ml_ms_n_24);
  ml_ms_g1896 : AOI22D0BWP7T port map(A1 => ml_ms_n_4, A2 => ml_ms_sr_new_new_data(7), B1 => ml_ms_n_9, B2 => ml_ms_sr_new_new_data(6), ZN => ml_ms_n_23);
  ml_ms_g1897 : AOI22D0BWP7T port map(A1 => ml_ms_n_4, A2 => ml_ms_sr_new_new_data(5), B1 => ml_ms_n_9, B2 => ml_ms_sr_new_new_data(4), ZN => ml_ms_n_22);
  ml_ms_g1898 : AOI22D0BWP7T port map(A1 => ml_ms_n_4, A2 => ml_ms_muxReg, B1 => ml_ms_n_9, B2 => ml_ms_sr_new_new_data(7), ZN => ml_ms_n_21);
  ml_ms_g1899 : AO22D0BWP7T port map(A1 => ml_ms_n_4, A2 => ml_ms_sr_new_new_data(1), B1 => ml_ms_sr_new_new_data(0), B2 => ml_ms_n_9, Z => FE_PHN459_ml_ms_n_20);
  ml_ms_g1900 : AO22D0BWP7T port map(A1 => ml_ms_n_4, A2 => ml_ms_sr_new_new_data(2), B1 => ml_ms_sr_new_new_data(1), B2 => ml_ms_n_9, Z => FE_PHN457_ml_ms_n_19);
  ml_ms_g1901 : INR2D1BWP7T port map(A1 => ml_ms_n_11, B1 => ml_ms_count25M(12), ZN => ml_ms_n_18);
  ml_ms_g1902 : INR2D1BWP7T port map(A1 => ml_ms_count25M(8), B1 => ml_ms_n_6, ZN => ml_ms_n_17);
  ml_ms_g1903 : OR2D1BWP7T port map(A1 => ml_ms_n_10, A2 => ml_ms_muxFSM, Z => ml_ms_n_16);
  ml_ms_g1904 : AOI21D0BWP7T port map(A1 => ml_ms_n_0, A2 => FE_PHN425_ml_ms_mux_select, B => ml_ms_muxFSM, ZN => ml_ms_n_14);
  ml_ms_g1905 : NR3D0BWP7T port map(A1 => ml_ms_count25M(3), A2 => FE_PHN437_ml_ms_count25M_4, A3 => ml_ms_count25M(5), ZN => ml_ms_n_13);
  ml_ms_g1906 : IAO21D0BWP7T port map(A1 => ml_ms_count25M(7), A2 => FE_PHN415_ml_ms_count25M_6, B => ml_ms_n_11, ZN => ml_ms_n_12);
  ml_ms_g1907 : NR3D0BWP7T port map(A1 => ml_ms_count25M(8), A2 => ml_ms_count25M(12), A3 => ml_ms_count25M(9), ZN => ml_ms_n_15);
  ml_ms_g1908 : ND2D1BWP7T port map(A1 => ml_ms_count25M(10), A2 => ml_ms_count25M(11), ZN => ml_ms_n_11);
  ml_ms_g1909 : IND2D1BWP7T port map(A1 => ml_ms_reset_send, B1 => FE_PHN416_ml_ms_sfsm_state_0, ZN => ml_ms_n_10);
  ml_ms_g1910 : AN2D1BWP7T port map(A1 => ml_ms_output_edgedet, A2 => FE_PHN425_ml_ms_mux_select, Z => ml_ms_n_9);
  ml_ms_g1911 : INVD1BWP7T port map(I => ml_ms_n_7, ZN => ml_ms_n_8);
  ml_ms_g1912 : INVD0BWP7T port map(I => ml_ms_n_6, ZN => ml_ms_n_5);
  ml_ms_g1913 : OR2D1BWP7T port map(A1 => FE_PHN437_ml_ms_count25M_4, A2 => ml_ms_count25M(2), Z => ml_ms_n_3);
  ml_ms_g1914 : NR2XD0BWP7T port map(A1 => ml_ms_reset_send, A2 => FE_PHN416_ml_ms_sfsm_state_0, ZN => ml_ms_n_7);
  ml_ms_g1915 : CKND2D1BWP7T port map(A1 => ml_ms_count25M(7), A2 => FE_PHN415_ml_ms_count25M_6, ZN => ml_ms_n_6);
  ml_ms_g1916 : NR2XD0BWP7T port map(A1 => ml_ms_output_edgedet, A2 => ml_ms_n_2, ZN => ml_ms_n_4);
  ml_ms_sfsm_state_reg_1 : DFD1BWP7T port map(CP => CTS_322, D => FE_PHN471_ml_ms_n_57, Q => ml_ms_sfsm_state(1), QN => ml_ms_n_0);
  ml_ms_sfsm_state_reg_3 : DFD1BWP7T port map(CP => CTS_288, D => FE_PHN469_ml_ms_n_60, Q => ml_ms_mux_select, QN => ml_ms_n_2);
  ml_ms_sfsm_state_reg_2 : DFD1BWP7T port map(CP => CTS_288, D => FE_PHN470_ml_ms_n_54, Q => ml_ms_muxFSM, QN => ml_ms_n_1);
  ml_ms_mfsm_g2084 : OR4D1BWP7T port map(A1 => ml_ms_mfsm_n_108, A2 => ml_ms_mfsm_n_110, A3 => ml_ms_mfsm_n_51, A4 => ml_ms_mfsm_n_57, Z => ml_ms_cntReset15K);
  ml_ms_mfsm_g2085 : AN2D0BWP7T port map(A1 => ml_ms_btnflipfloprst, A2 => ml_ms_data_sr_11bit(3), Z => ml_ms_btns(4));
  ml_ms_mfsm_g2086 : AN2D0BWP7T port map(A1 => ml_ms_btnflipfloprst, A2 => ml_ms_data_sr_11bit(4), Z => ml_ms_btns(3));
  ml_ms_mfsm_g2087 : AN2D0BWP7T port map(A1 => ml_ms_btnflipfloprst, A2 => ml_ms_data_sr_11bit(2), Z => ml_ms_btns(2));
  ml_ms_mfsm_g2088 : AN2D0BWP7T port map(A1 => ml_ms_btnflipfloprst, A2 => FE_PHN411_ml_ms_data_sr_11bit_7, Z => ml_ms_btns(1));
  ml_ms_mfsm_g2089 : AN2D0BWP7T port map(A1 => ml_ms_btnflipfloprst, A2 => ml_ms_data_sr_11bit(6), Z => ml_ms_btns(0));
  ml_ms_mfsm_g2090 : INR2D1BWP7T port map(A1 => ml_ms_data_sr_11bit(2), B1 => ml_ms_mfsm_n_58, ZN => ml_ms_mouse_x(0));
  ml_ms_mfsm_g2091 : INR2D1BWP7T port map(A1 => ml_ms_data_sr_11bit(3), B1 => ml_ms_mfsm_n_58, ZN => ml_ms_mouse_x(1));
  ml_ms_mfsm_g2092 : INR2D1BWP7T port map(A1 => ml_ms_data_sr_11bit(4), B1 => ml_ms_mfsm_n_58, ZN => ml_ms_mouse_x(2));
  ml_ms_mfsm_g2093 : AN2D0BWP7T port map(A1 => ml_ms_yflipfloprst, A2 => ml_ms_data_sr_11bit(4), Z => ml_ms_mouse_y(2));
  ml_ms_mfsm_g2094 : AN2D0BWP7T port map(A1 => ml_ms_yflipfloprst, A2 => ml_ms_data_sr_11bit(2), Z => ml_ms_mouse_y(0));
  ml_ms_mfsm_g2095 : AN2D0BWP7T port map(A1 => ml_ms_yflipfloprst, A2 => ml_ms_data_sr_11bit(3), Z => ml_ms_mouse_y(1));
  ml_ms_mfsm_g2096 : ND3D0BWP7T port map(A1 => ml_ms_mfsm_n_54, A2 => ml_ms_mfsm_n_55, A3 => ml_ms_mfsm_state(1), ZN => ml_ms_cntReset25M_main);
  ml_ms_mfsm_g2097 : OAI31D1BWP7T port map(A1 => ml_ms_mfsm_state(3), A2 => ml_ms_mfsm_state(2), A3 => ml_ms_mfsm_n_52, B => ml_ms_mfsm_n_56, ZN => FE_PHN486_ml_ms_btnflipfloprst);
  ml_ms_mfsm_g2098 : IAO21D0BWP7T port map(A1 => ml_ms_mfsm_n_52, A2 => ml_ms_mfsm_n_47, B => ml_ms_xflipfloprst, ZN => ml_ms_mfsm_n_58);
  ml_ms_mfsm_g2099 : OAI21D0BWP7T port map(A1 => ml_ms_mfsm_n_53, A2 => FE_PHN454_ml_ms_mfsm_state_0, B => ml_ms_mfsm_n_56, ZN => ml_ms_mfsm_n_57);
  ml_ms_mfsm_g2100 : MOAI22D0BWP7T port map(A1 => ml_ms_mfsm_n_52, A2 => ml_ms_mfsm_n_0, B1 => ml_ms_mfsm_n_110, B2 => ml_ms_mfsm_state(2), ZN => ml_ms_yflipfloprst);
  ml_ms_mfsm_g2101 : IND2D1BWP7T port map(A1 => ml_ms_mfsm_n_51, B1 => ml_ms_mfsm_n_53, ZN => ml_ms_mux_select_main);
  ml_ms_mfsm_g2102 : NR2XD0BWP7T port map(A1 => ml_ms_reset_send, A2 => ml_ms_mfsm_n_0, ZN => ml_ms_actBit);
  ml_ms_mfsm_g2103 : AN2D1BWP7T port map(A1 => ml_ms_mfsm_n_110, A2 => ml_ms_mfsm_n_47, Z => ml_ms_xflipfloprst);
  ml_ms_mfsm_g2104 : AOI22D0BWP7T port map(A1 => ml_ms_mfsm_n_50, A2 => ml_ms_mfsm_state(2), B1 => ml_ms_mfsm_n_47, B2 => ml_ms_mfsm_state(3), ZN => ml_ms_mfsm_n_55);
  ml_ms_mfsm_g2105 : MAOI22D0BWP7T port map(A1 => ml_ms_mfsm_n_48, A2 => FE_PHN454_ml_ms_mfsm_state_0, B1 => ml_ms_mfsm_n_48, B2 => FE_PHN454_ml_ms_mfsm_state_0, ZN => ml_ms_mfsm_n_54);
  ml_ms_mfsm_g2106 : ND3D0BWP7T port map(A1 => ml_ms_mfsm_n_60, A2 => ml_ms_mfsm_state(2), A3 => ml_ms_mfsm_state(3), ZN => ml_ms_mfsm_n_56);
  ml_ms_mfsm_g2107 : INR2D1BWP7T port map(A1 => ml_ms_mfsm_n_48, B1 => ml_ms_mfsm_n_50, ZN => ml_ms_mfsm_n_53);
  ml_ms_mfsm_g2108 : ND2D1BWP7T port map(A1 => ml_ms_mfsm_n_49, A2 => ml_ms_mfsm_state(4), ZN => ml_ms_mfsm_n_52);
  ml_ms_mfsm_g2109 : AN2D1BWP7T port map(A1 => ml_ms_mfsm_n_60, A2 => ml_ms_mfsm_state(4), Z => ml_ms_mfsm_n_110);
  ml_ms_mfsm_g2110 : AN2D0BWP7T port map(A1 => ml_ms_mfsm_n_108, A2 => FE_PHN454_ml_ms_mfsm_state_0, Z => ml_handshake_mouse_out);
  ml_ms_mfsm_g2111 : IND2D1BWP7T port map(A1 => ml_ms_mfsm_n_48, B1 => ml_ms_mfsm_n_109, ZN => ml_ms_reset_send);
  ml_ms_mfsm_g2112 : CKAN2D1BWP7T port map(A1 => ml_ms_mfsm_n_49, A2 => ml_ms_mfsm_n_2, Z => ml_ms_mfsm_n_51);
  ml_ms_mfsm_g2113 : INR2XD0BWP7T port map(A1 => FE_PHN454_ml_ms_mfsm_state_0, B1 => ml_ms_mfsm_state(1), ZN => ml_ms_mfsm_n_109);
  ml_ms_mfsm_g2114 : AN2D1BWP7T port map(A1 => ml_ms_mfsm_state(1), A2 => FE_PHN454_ml_ms_mfsm_state_0, Z => ml_ms_mfsm_n_60);
  ml_ms_mfsm_g2115 : NR2D1BWP7T port map(A1 => ml_ms_mfsm_n_2, A2 => ml_ms_mfsm_n_0, ZN => ml_ms_mfsm_n_108);
  ml_ms_mfsm_g2116 : ND2D1BWP7T port map(A1 => ml_ms_mfsm_state(4), A2 => FE_PHN454_ml_ms_mfsm_state_0, ZN => ml_ms_mfsm_n_57_BAR);
  ml_ms_mfsm_g2117 : NR2XD0BWP7T port map(A1 => ml_ms_mfsm_state(4), A2 => ml_ms_mfsm_state(3), ZN => ml_ms_mfsm_n_50);
  ml_ms_mfsm_g2118 : NR2XD0BWP7T port map(A1 => ml_ms_mfsm_state(1), A2 => FE_PHN454_ml_ms_mfsm_state_0, ZN => ml_ms_mfsm_n_49);
  ml_ms_mfsm_g2119 : ND2D1BWP7T port map(A1 => ml_ms_mfsm_n_2, A2 => ml_ms_mfsm_n_47, ZN => ml_ms_mfsm_n_48);
  ml_ms_mfsm_state_reg_0 : DFQD1BWP7T port map(CP => CTS_322, D => ml_ms_mfsm_n_46, Q => ml_ms_mfsm_state(0));
  ml_ms_mfsm_state_reg_1 : DFQD1BWP7T port map(CP => CTS_322, D => FE_PHN477_ml_ms_mfsm_n_45, Q => ml_ms_mfsm_state(1));
  ml_ms_mfsm_g2643 : OAI31D0BWP7T port map(A1 => FE_OFN31_reset, A2 => ml_ms_mfsm_n_21, A3 => ml_ms_mfsm_n_30, B => ml_ms_mfsm_n_44, ZN => FE_PHN478_ml_ms_mfsm_n_46);
  ml_ms_mfsm_g2644 : AO222D0BWP7T port map(A1 => ml_ms_mfsm_n_40, A2 => ml_ms_mfsm_state(1), B1 => ml_handshake_mouse_out, B2 => ml_ms_mfsm_n_7, C1 => ml_ms_mfsm_n_37, C2 => FE_PHN454_ml_ms_mfsm_state_0, Z => ml_ms_mfsm_n_45);
  ml_ms_mfsm_g2645 : AOI211XD0BWP7T port map(A1 => ml_ms_mfsm_n_19, A2 => ml_ms_count25M(12), B => ml_ms_mfsm_n_41, C => ml_ms_mfsm_n_20, ZN => ml_ms_mfsm_n_44);
  ml_ms_mfsm_g2648 : OAI211D1BWP7T port map(A1 => ml_ms_mfsm_state(4), A2 => ml_ms_mfsm_n_33, B => ml_ms_mfsm_n_39, C => ml_ms_mfsm_n_16, ZN => ml_ms_mfsm_n_43);
  ml_ms_mfsm_g2649 : OAI32D1BWP7T port map(A1 => ml_ms_mfsm_state(3), A2 => ml_ms_mfsm_n_6, A3 => ml_ms_mfsm_n_35, B1 => FE_OFN31_reset, B2 => ml_ms_mfsm_n_26, ZN => FE_PHN466_ml_ms_mfsm_n_42);
  ml_ms_mfsm_g2650 : MOAI22D0BWP7T port map(A1 => ml_ms_mfsm_n_38, A2 => ml_ms_mfsm_n_18, B1 => ml_ms_mfsm_n_31, B2 => ml_ms_mfsm_n_27, ZN => ml_ms_mfsm_n_41);
  ml_ms_mfsm_g2651 : OAI221D0BWP7T port map(A1 => ml_ms_mfsm_n_32, A2 => ml_ms_mfsm_state(4), B1 => ml_ms_mfsm_state(4), B2 => ml_ms_mfsm_n_33, C => ml_ms_mfsm_n_18, ZN => ml_ms_mfsm_n_40);
  ml_ms_mfsm_g2652 : AOI32D1BWP7T port map(A1 => ml_ms_mfsm_n_10, A2 => ml_ms_mfsm_state(4), A3 => ml_ms_mfsm_n_11, B1 => ml_ms_mfsm_n_36, B2 => ml_ms_mfsm_n_8, ZN => ml_ms_mfsm_n_39);
  ml_ms_mfsm_g2653 : OAI31D0BWP7T port map(A1 => ml_ms_count25M(9), A2 => ml_ms_count25M(10), A3 => ml_ms_mfsm_n_28, B => ml_ms_count25M(11), ZN => ml_ms_mfsm_n_38);
  ml_ms_mfsm_g2654 : MOAI22D0BWP7T port map(A1 => ml_ms_mfsm_n_34, A2 => ml_ms_mfsm_state(1), B1 => ml_ms_mfsm_n_10, B2 => ml_ms_mfsm_n_12, ZN => ml_ms_mfsm_n_37);
  ml_ms_mfsm_g2655 : INVD0BWP7T port map(I => ml_ms_mfsm_n_35, ZN => ml_ms_mfsm_n_36);
  ml_ms_mfsm_g2656 : AOI21D0BWP7T port map(A1 => ml_ms_mfsm_n_30, A2 => ml_ms_mfsm_state(1), B => ml_ms_mfsm_n_110, ZN => ml_ms_mfsm_n_35);
  ml_ms_mfsm_g2657 : OAI21D0BWP7T port map(A1 => ml_ms_mfsm_n_22, A2 => ml_ms_mfsm_n_5, B => FE_PHN417_ml_ms_count15k_3, ZN => ml_ms_mfsm_n_34);
  ml_ms_mfsm_g2659 : AOI21D0BWP7T port map(A1 => ml_ms_mfsm_n_23, A2 => ml_ms_mfsm_n_8, B => ml_ms_mfsm_n_11, ZN => ml_ms_mfsm_n_32);
  ml_ms_mfsm_g2660 : OAI21D0BWP7T port map(A1 => FE_PHN422_ml_ms_count15k_2, A2 => ml_ms_mfsm_state(1), B => ml_ms_mfsm_n_30, ZN => ml_ms_mfsm_n_31);
  ml_ms_mfsm_g2661 : ND3D0BWP7T port map(A1 => ml_ms_mfsm_n_23, A2 => ml_ms_mfsm_n_7, A3 => ml_ms_mfsm_n_0, ZN => ml_ms_mfsm_n_33);
  ml_ms_mfsm_g2662 : OAI211D1BWP7T port map(A1 => FE_OFN31_reset, A2 => ml_ms_mfsm_n_57_BAR, B => ml_ms_mfsm_n_25, C => ml_ms_mfsm_n_17, ZN => FE_PHN473_ml_ms_mfsm_n_29);
  ml_ms_mfsm_g2663 : INR2XD0BWP7T port map(A1 => FE_PHN454_ml_ms_mfsm_state_0, B1 => ml_ms_mfsm_n_23, ZN => ml_ms_mfsm_n_30);
  ml_ms_mfsm_g2664 : AN4D0BWP7T port map(A1 => ml_ms_mfsm_n_15, A2 => FE_PHN415_ml_ms_count25M_6, A3 => ml_ms_count25M(7), A4 => ml_ms_count25M(8), Z => ml_ms_mfsm_n_28);
  ml_ms_mfsm_g2665 : AO21D0BWP7T port map(A1 => ml_ms_mfsm_n_8, A2 => ml_ms_mfsm_n_2, B => ml_ms_mfsm_n_24, Z => ml_ms_mfsm_n_27);
  ml_ms_mfsm_g2666 : AOI21D0BWP7T port map(A1 => ml_ms_mfsm_n_4, A2 => ml_ms_mfsm_state(3), B => ml_ms_mfsm_n_10, ZN => ml_ms_mfsm_n_26);
  ml_ms_mfsm_g2667 : OAI211D1BWP7T port map(A1 => ml_ms_mfsm_state(4), A2 => ml_ms_mfsm_n_60, B => ml_ms_mfsm_n_7, C => ml_ms_mfsm_state(3), ZN => ml_ms_mfsm_n_25);
  ml_ms_mfsm_g2668 : NR3D0BWP7T port map(A1 => ml_ms_mfsm_n_109, A2 => ml_ms_mfsm_n_9, A3 => FE_OFN31_reset, ZN => ml_ms_mfsm_n_24);
  ml_ms_mfsm_g2669 : IAO21D0BWP7T port map(A1 => ml_ms_mfsm_n_7, A2 => ml_ms_mfsm_n_12, B => ml_ms_tb_n_2, ZN => ml_ms_mfsm_n_22);
  ml_ms_mfsm_g2670 : OA22D0BWP7T port map(A1 => ml_ms_mfsm_n_10, A2 => ml_ms_mfsm_state(1), B1 => ml_ms_mfsm_state(4), B2 => ml_ms_mfsm_state(3), Z => ml_ms_mfsm_n_21);
  ml_ms_mfsm_g2671 : NR4D0BWP7T port map(A1 => ml_ms_mfsm_n_6, A2 => ml_ms_mfsm_n_0, A3 => ml_ms_mfsm_state(4), A4 => ml_ms_mfsm_state(1), ZN => ml_ms_mfsm_n_20);
  ml_ms_mfsm_g2672 : OAI21D0BWP7T port map(A1 => ml_ms_mfsm_n_14, A2 => FE_PHN422_ml_ms_count15k_2, B => FE_PHN417_ml_ms_count15k_3, ZN => ml_ms_mfsm_n_23);
  ml_ms_mfsm_g2673 : INVD0BWP7T port map(I => ml_ms_mfsm_n_18, ZN => ml_ms_mfsm_n_19);
  ml_ms_mfsm_g2674 : ND2D1BWP7T port map(A1 => ml_ms_mfsm_n_12, A2 => ml_ms_mfsm_n_0, ZN => ml_ms_mfsm_n_17);
  ml_ms_mfsm_g2675 : ND2D1BWP7T port map(A1 => ml_ms_mfsm_n_9, A2 => ml_ms_mfsm_n_11, ZN => ml_ms_mfsm_n_18);
  ml_ms_mfsm_g2676 : OAI21D0BWP7T port map(A1 => ml_ms_mfsm_n_1, A2 => ml_ms_mfsm_n_108, B => ml_ms_mfsm_n_7, ZN => ml_ms_mfsm_n_16);
  ml_ms_mfsm_g2677 : OR4D1BWP7T port map(A1 => ml_ms_count25M(5), A2 => FE_PHN437_ml_ms_count25M_4, A3 => ml_ms_count25M(3), A4 => ml_ms_count25M(2), Z => ml_ms_mfsm_n_15);
  ml_ms_mfsm_g2678 : INVD1BWP7T port map(I => ml_ms_tb_n_2, ZN => ml_ms_mfsm_n_14);
  ml_ms_mfsm_g2679 : INVD0BWP7T port map(I => ml_ms_mfsm_n_10, ZN => ml_ms_mfsm_n_9);
  ml_ms_mfsm_g2681 : NR2D1BWP7T port map(A1 => ml_ms_mfsm_n_2, A2 => FE_OFN31_reset, ZN => ml_ms_mfsm_n_12);
  ml_ms_mfsm_g2682 : NR2D1BWP7T port map(A1 => FE_PHN454_ml_ms_mfsm_state_0, A2 => FE_OFN31_reset, ZN => ml_ms_mfsm_n_11);
  ml_ms_mfsm_g2683 : NR2D1BWP7T port map(A1 => ml_ms_mfsm_n_0, A2 => ml_ms_mfsm_state(2), ZN => ml_ms_mfsm_n_10);
  ml_ms_mfsm_g2684 : INVD0BWP7T port map(I => ml_ms_mfsm_n_7, ZN => ml_ms_mfsm_n_6);
  ml_ms_mfsm_g2685 : INR2D1BWP7T port map(A1 => FE_PHN422_ml_ms_count15k_2, B1 => FE_OFN31_reset, ZN => ml_ms_mfsm_n_5);
  ml_ms_mfsm_g2686 : ND2D1BWP7T port map(A1 => ml_ms_mfsm_n_60, A2 => ml_ms_mfsm_n_2, ZN => ml_ms_mfsm_n_4);
  ml_ms_mfsm_g2687 : NR2XD0BWP7T port map(A1 => ml_ms_mfsm_state(2), A2 => FE_OFN31_reset, ZN => ml_ms_mfsm_n_8);
  ml_ms_mfsm_g2688 : INR2D1BWP7T port map(A1 => ml_ms_mfsm_state(2), B1 => FE_OFN31_reset, ZN => ml_ms_mfsm_n_7);
  ml_ms_mfsm_g2691 : INVD0BWP7T port map(I => ml_ms_mfsm_n_60, ZN => ml_ms_mfsm_n_1);
  ml_ms_mfsm_state_reg_4 : DFD1BWP7T port map(CP => CTS_322, D => ml_ms_mfsm_n_29, Q => ml_ms_mfsm_state(4), QN => ml_ms_mfsm_n_2);
  ml_ms_mfsm_state_reg_3 : DFD1BWP7T port map(CP => CTS_322, D => ml_ms_mfsm_n_42, Q => ml_ms_mfsm_state(3), QN => ml_ms_mfsm_n_0);
  ml_ms_mfsm_state_reg_2 : DFD1BWP7T port map(CP => CTS_322, D => FE_PHN476_ml_ms_mfsm_n_43, Q => FE_PHN443_ml_ms_mfsm_state_2, QN => FE_PHN452_ml_ms_mfsm_n_47);
  ml_ms_flipflop10_Q_reg : DFXQD1BWP7T port map(CP => CTS_322, DA => ml_ms_btns(1), DB => FE_PHN420_ml_buttons_mouse_1, Q => ml_buttons_mouse(1), SA => ml_ms_btnflipfloprst);
  ml_ms_flipflop1_Q_reg : DFXQD1BWP7T port map(CP => CTS_322, DA => ml_ms_mouse_x(2), DB => ml_mouseX(2), Q => FE_PHN429_ml_mouseX_2, SA => ml_ms_xflipfloprst);
  ml_ms_tb_count_reg_3 : EDFKCNQD1BWP7T port map(CN => ml_ms_tb_n_1, CP => CTS_322, D => ml_ms_tb_n_6, E => ml_ms_output_edgedet, Q => ml_ms_count15k(3));
  ml_ms_tb_count_reg_2 : EDFKCNQD1BWP7T port map(CN => ml_ms_tb_n_1, CP => CTS_322, D => FE_PHN509_ml_ms_tb_n_5, E => ml_ms_output_edgedet, Q => ml_ms_count15k(2));
  ml_ms_tb_g65 : MOAI22D0BWP7T port map(A1 => ml_ms_tb_n_4, A2 => FE_PHN417_ml_ms_count15k_3, B1 => ml_ms_tb_n_4, B2 => FE_PHN417_ml_ms_count15k_3, ZN => FE_PHN475_ml_ms_tb_n_6);
  ml_ms_tb_count_reg_1 : EDFKCNQD1BWP7T port map(CN => ml_ms_tb_n_1, CP => CTS_322, D => ml_ms_tb_n_3, E => ml_ms_output_edgedet, Q => FE_PHN504_ml_ms_count15k_1);
  ml_ms_tb_g67 : MOAI22D0BWP7T port map(A1 => ml_ms_tb_n_2, A2 => FE_PHN422_ml_ms_count15k_2, B1 => ml_ms_tb_n_2, B2 => FE_PHN422_ml_ms_count15k_2, ZN => ml_ms_tb_n_5);
  ml_ms_tb_count_reg_0 : DFKCNQD1BWP7T port map(CN => ml_ms_tb_n_0, CP => CTS_322, D => ml_ms_tb_n_1, Q => FE_PHN414_ml_ms_count15k_0);
  ml_ms_tb_g69 : IND2D1BWP7T port map(A1 => ml_ms_tb_n_2, B1 => FE_PHN422_ml_ms_count15k_2, ZN => ml_ms_tb_n_4);
  ml_ms_tb_g70 : CKXOR2D0BWP7T port map(A1 => ml_ms_count15k(1), A2 => ml_ms_count15k(0), Z => ml_ms_tb_n_3);
  ml_ms_tb_g72 : ND2D1BWP7T port map(A1 => ml_ms_count15k(1), A2 => ml_ms_count15k(0), ZN => ml_ms_tb_n_2);
  ml_ms_tb_g73 : INVD1BWP7T port map(I => ml_ms_cntReset15K, ZN => ml_ms_tb_n_1);
  ml_ms_tb_g2 : CKXOR2D1BWP7T port map(A1 => ml_ms_output_edgedet, A2 => ml_ms_count15k(0), Z => ml_ms_tb_n_0);
  ml_ms_flipflop11_Q_reg : DFXQD1BWP7T port map(CP => CTS_322, DA => ml_ms_btns(0), DB => ml_buttons_mouse(0), Q => FE_PHN440_ml_buttons_mouse_0, SA => ml_ms_btnflipfloprst);
  ml_ms_flipflop2_Q_reg : DFXQD1BWP7T port map(CP => CTS_322, DA => ml_ms_mouse_x(1), DB => FE_PHN391_ml_mouseX_1, Q => ml_mouseX(1), SA => ml_ms_xflipfloprst);
  ml_ms_sr11_data_out_reg_1 : EDFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_288, D => FE_PHN387_ml_ms_sr11_data_out_0_79, E => ml_ms_output_edgedet, Q => ml_ms_sr11_data_out_1_80);
  ml_ms_sr11_data_out_reg_0 : EDFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_288, D => FE_PHN404_data_in, E => ml_ms_output_edgedet, Q => ml_ms_sr11_data_out_0_79);
  ml_ms_sr11_data_out_reg_3 : EDFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_322, D => ml_ms_data_sr_11bit(2), E => ml_ms_output_edgedet, Q => FE_PHN380_ml_ms_data_sr_11bit_3);
  ml_ms_sr11_data_out_reg_4 : EDFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_322, D => ml_ms_data_sr_11bit(3), E => ml_ms_output_edgedet, Q => FE_PHN385_ml_ms_data_sr_11bit_4);
  ml_ms_sr11_data_out_reg_5 : EDFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_322, D => ml_ms_data_sr_11bit(4), E => ml_ms_output_edgedet, Q => FE_PHN388_ml_ms_sr11_data_out_5_84);
  ml_ms_sr11_data_out_reg_7 : EDFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_322, D => ml_ms_data_sr_11bit(6), E => ml_ms_output_edgedet, Q => ml_ms_data_sr_11bit(7));
  ml_ms_sr11_data_out_reg_6 : EDFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_322, D => ml_ms_sr11_data_out_5_84, E => ml_ms_output_edgedet, Q => FE_PHN383_ml_ms_data_sr_11bit_6);
  ml_ms_sr11_data_out_reg_2 : EDFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_288, D => FE_PHN390_ml_ms_sr11_data_out_1_80, E => ml_ms_output_edgedet, Q => FE_PHN386_ml_ms_data_sr_11bit_2);
  ml_ms_flipflop3_Q_reg : DFXQD1BWP7T port map(CP => CTS_322, DA => ml_ms_mouse_x(0), DB => FE_PHN398_ml_mouseX_0, Q => ml_mouseX(0), SA => ml_ms_xflipfloprst);
  ml_ms_flipflop4_Q_reg : DFXQD1BWP7T port map(CP => CTS_322, DA => ml_ms_mouse_y(0), DB => FE_PHN401_ml_mouseY_0, Q => ml_mouseY(0), SA => ml_ms_yflipfloprst);
  ml_il_y1_g531 : OAI222D0BWP7T port map(A1 => ml_il_y1_n_27, A2 => ml_il_y1_n_6, B1 => ml_il_y1_n_3, B2 => ml_il_y1_cmbsop_sel(1), C1 => ml_il_y1_n_8, C2 => ml_il_y1_n_29, ZN => ml_il_y1_input_register(3));
  ml_il_y1_g532 : MAOI22D0BWP7T port map(A1 => ml_il_y1_n_28, A2 => ml_il_y1_input_register(3), B1 => ml_il_y1_n_28, B2 => ml_il_y1_input_register(3), ZN => ml_il_y1_n_29);
  ml_il_y1_g533 : AO21D0BWP7T port map(A1 => ml_il_y1_n_25, A2 => ml_il_y1_n_17, B => ml_il_y1_n_20, Z => ml_il_y1_n_28);
  ml_il_y1_g534 : MAOI22D0BWP7T port map(A1 => ml_il_y1_n_26, A2 => ml_il_y1_input_register(3), B1 => ml_il_y1_n_26, B2 => ml_il_y1_input_register(3), ZN => ml_il_y1_n_27);
  ml_il_y1_g535 : MOAI22D0BWP7T port map(A1 => ml_il_y1_n_25, A2 => ml_il_y1_n_23, B1 => ml_il_y1_n_25, B2 => ml_il_y1_n_23, ZN => ml_il_y1_n_40);
  ml_il_y1_g536 : MAOI222D1BWP7T port map(A => ml_il_y1_n_24, B => ml_il_y1_n_49, C => FE_PHN392_ml_mouseY_2, ZN => ml_il_y1_n_26);
  ml_il_y1_g537 : AO21D0BWP7T port map(A1 => ml_il_y1_n_16, A2 => ml_il_y1_n_21, B => ml_il_y1_n_18, Z => ml_il_y1_n_25);
  ml_il_y1_g538 : CKXOR2D0BWP7T port map(A1 => ml_il_y1_n_24, A2 => ml_il_y1_n_23, Z => ml_il_y1_n_39);
  ml_il_y1_g539 : MOAI22D0BWP7T port map(A1 => ml_il_y1_n_22, A2 => ml_il_y1_n_16, B1 => ml_il_y1_n_22, B2 => ml_il_y1_n_16, ZN => ml_il_y1_n_42);
  ml_il_y1_g540 : MOAI22D0BWP7T port map(A1 => ml_il_y1_n_22, A2 => ml_il_y1_n_19, B1 => ml_il_y1_n_22, B2 => ml_il_y1_n_19, ZN => ml_il_y1_n_41);
  ml_il_y1_g541 : MAOI222D1BWP7T port map(A => ml_il_y1_n_19, B => ml_il_y1_n_14, C => ml_il_y1_n_4, ZN => ml_il_y1_n_24);
  ml_il_y1_g542 : IND2D0BWP7T port map(A1 => ml_il_y1_n_20, B1 => ml_il_y1_n_17, ZN => ml_il_y1_n_23);
  ml_il_y1_g543 : OAI21D0BWP7T port map(A1 => ml_il_y1_n_15, A2 => ml_mouseY(0), B => ml_il_y1_n_16, ZN => ml_il_y1_n_43);
  ml_il_y1_g544 : IND2D0BWP7T port map(A1 => ml_il_y1_n_18, B1 => ml_il_y1_n_21, ZN => ml_il_y1_n_22);
  ml_il_y1_g545 : ND2D1BWP7T port map(A1 => ml_il_y1_n_14, A2 => FE_PHN395_ml_mouseY_1, ZN => ml_il_y1_n_21);
  ml_il_y1_g546 : NR2D0BWP7T port map(A1 => ml_il_y1_n_13, A2 => FE_PHN392_ml_mouseY_2, ZN => ml_il_y1_n_20);
  ml_il_y1_g547 : ND2D1BWP7T port map(A1 => ml_il_y1_n_47, A2 => ml_mouseY(0), ZN => ml_il_y1_n_19);
  ml_il_y1_g548 : NR2D0BWP7T port map(A1 => ml_il_y1_n_14, A2 => FE_PHN395_ml_mouseY_1, ZN => ml_il_y1_n_18);
  ml_il_y1_g549 : ND2D1BWP7T port map(A1 => ml_il_y1_n_13, A2 => FE_PHN392_ml_mouseY_2, ZN => ml_il_y1_n_17);
  ml_il_y1_g550 : ND2D1BWP7T port map(A1 => ml_il_y1_n_15, A2 => ml_mouseY(0), ZN => ml_il_y1_n_16);
  ml_il_y1_g551 : CKND1BWP7T port map(I => ml_il_y1_n_47, ZN => ml_il_y1_n_15);
  ml_il_y1_g553 : INVD1BWP7T port map(I => ml_il_y1_n_48, ZN => ml_il_y1_n_14);
  ml_il_y1_g554 : CKND1BWP7T port map(I => ml_il_y1_n_49, ZN => ml_il_y1_n_13);
  ml_il_y1_g560 : INVD1BWP7T port map(I => ml_il_y1_n_8, ZN => ml_il_y1_n_9);
  ml_il_y1_g561 : ND2D1BWP7T port map(A1 => ml_il_y1_cmbsop_sel(1), A2 => FE_PHN420_ml_buttons_mouse_1, ZN => ml_il_y1_n_8);
  ml_il_y1_g562 : INVD0BWP7T port map(I => ml_il_y1_n_7, ZN => ml_il_y1_n_6);
  ml_il_y1_g563 : NR2XD0BWP7T port map(A1 => ml_il_y1_n_5, A2 => FE_PHN420_ml_buttons_mouse_1, ZN => ml_il_y1_n_7);
  ml_il_y1_g564 : INVD1BWP7T port map(I => ml_il_y1_cmbsop_sel(1), ZN => ml_il_y1_n_5);
  ml_il_y1_g565 : INR2D1BWP7T port map(A1 => FE_PHN424_ml_il_y1_state_0, B1 => FE_PHN402_ml_il_y1_state_1, ZN => ml_il_y1_cmbsop_sel(1));
  ml_il_y1_g566 : INVD0BWP7T port map(I => FE_PHN395_ml_mouseY_1, ZN => ml_il_y1_n_4);
  ml_il_y1_state_reg_0 : DFQD1BWP7T port map(CP => CTS_322, D => ml_il_y1_n_2, Q => ml_il_y1_state(0));
  ml_il_y1_state_reg_1 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_322, D => ml_il_y1_n_1, Q => ml_il_y1_state(1));
  ml_il_y1_g255 : INR4D0BWP7T port map(A1 => ml_handshake_mouse_out, B1 => FE_OFN31_reset, B2 => FE_PHN402_ml_il_y1_state_1, B3 => FE_PHN424_ml_il_y1_state_0, ZN => ml_il_y1_n_2);
  ml_il_y1_tempy_reg_0 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_322, D => FE_PHN485_ml_il_y1_n_47, Q => sig_logic_y(0));
  ml_il_y1_tempy_reg_1 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_322, D => FE_PHN482_ml_il_y1_n_48, Q => sig_logic_y(1));
  ml_il_y1_tempy_reg_2 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_322, D => FE_PHN479_ml_il_y1_n_49, Q => sig_logic_y(2));
  ml_il_y1_g260 : AO21D0BWP7T port map(A1 => ml_handshake_mouse_out, A2 => FE_PHN402_ml_il_y1_state_1, B => ml_il_y1_cmbsop_sel(1), Z => ml_il_y1_n_1);
  ml_il_y1_tempy_reg_3 : DFKCND1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_322, D => FE_PHN483_ml_il_y1_input_register_3, Q => sig_logic_y(3), QN => ml_il_y1_n_3);
  ml_il_y1_g2 : AO222D0BWP7T port map(A1 => ml_il_y1_n_7, A2 => ml_il_y1_n_43, B1 => ml_il_y1_n_9, B2 => ml_il_y1_n_43, C1 => ml_il_y1_n_5, C2 => sig_logic_y(0), Z => ml_il_y1_n_47);
  ml_il_y1_g570 : AO222D0BWP7T port map(A1 => ml_il_y1_n_7, A2 => ml_il_y1_n_41, B1 => ml_il_y1_n_9, B2 => ml_il_y1_n_42, C1 => ml_il_y1_n_5, C2 => sig_logic_y(1), Z => ml_il_y1_n_48);
  ml_il_y1_g571 : AO222D0BWP7T port map(A1 => ml_il_y1_n_7, A2 => ml_il_y1_n_39, B1 => ml_il_y1_n_9, B2 => ml_il_y1_n_40, C1 => ml_il_y1_n_5, C2 => FE_PHN530_sig_logic_y_2, Z => ml_il_y1_n_49);
  ml_ms_flipflop5_Q_reg : DFXQD1BWP7T port map(CP => CTS_322, DA => ml_ms_mouse_y(1), DB => FE_PHN395_ml_mouseY_1, Q => ml_mouseY(1), SA => ml_ms_yflipfloprst);
  ml_ms_flipflop6_Q_reg : DFXQD1BWP7T port map(CP => CTS_322, DA => ml_ms_mouse_y(2), DB => FE_PHN392_ml_mouseY_2, Q => ml_mouseY(2), SA => ml_ms_yflipfloprst);
  ml_ms_flipflop7_Q_reg : DFXQD1BWP7T port map(CP => CTS_322, DA => ml_ms_btns(4), DB => FE_PHN381_ml_buttons_mouse_4, Q => ml_buttons_mouse(4), SA => ml_ms_btnflipfloprst);
  ml_ms_flipflop8_Q_reg : DFXQD1BWP7T port map(CP => CTS_322, DA => ml_ms_btns(3), DB => FE_PHN358_ml_buttons_mouse_3, Q => ml_buttons_mouse(3), SA => ml_ms_btnflipfloprst);
  ml_ms_mx_g23 : ND2D5BWP7T port map(A1 => ml_ms_mx_n_0, A2 => ml_ms_mx_n_1, ZN => data_switch);
  ml_ms_mx_g24 : ND2D1BWP7T port map(A1 => FE_PHN425_ml_ms_mux_select, A2 => ml_ms_muxReg, ZN => ml_ms_mx_n_1);
  ml_ms_mx_g25 : IND2D1BWP7T port map(A1 => FE_PHN425_ml_ms_mux_select, B1 => ml_ms_muxFSM, ZN => ml_ms_mx_n_0);
  ml_ms_flipflop9_Q_reg : DFXQD1BWP7T port map(CP => CTS_288, DA => ml_ms_btns(2), DB => FE_PHN394_ml_buttons_mouse_2, Q => ml_buttons_mouse(2), SA => ml_ms_btnflipfloprst);
  ml_ms_cnt_g71 : CKND1BWP7T port map(I => ml_ms_cntReset25M, ZN => ml_ms_cnt_n_23);
  ml_ms_cnt_count_reg_12 : DFKCNQD1BWP7T port map(CN => ml_ms_cnt_n_23, CP => CTS_288, D => FE_PHN493_ml_ms_cnt_n_22, Q => ml_ms_count25M(12));
  ml_ms_cnt_count_reg_11 : DFKCNQD1BWP7T port map(CN => ml_ms_cnt_n_23, CP => CTS_288, D => ml_ms_cnt_n_21, Q => ml_ms_count25M(11));
  ml_ms_cnt_g225 : MOAI22D0BWP7T port map(A1 => ml_ms_cnt_n_20, A2 => ml_ms_count25M(12), B1 => ml_ms_cnt_n_20, B2 => ml_ms_count25M(12), ZN => ml_ms_cnt_n_22);
  ml_ms_cnt_count_reg_10 : DFKCNQD1BWP7T port map(CN => ml_ms_cnt_n_23, CP => CTS_288, D => FE_PHN492_ml_ms_cnt_n_19, Q => FE_PHN427_ml_ms_count25M_10);
  ml_ms_cnt_g227 : MOAI22D0BWP7T port map(A1 => ml_ms_cnt_n_18, A2 => ml_ms_count25M(11), B1 => ml_ms_cnt_n_18, B2 => ml_ms_count25M(11), ZN => FE_PHN494_ml_ms_cnt_n_21);
  ml_ms_cnt_g228 : IND2D1BWP7T port map(A1 => ml_ms_cnt_n_18, B1 => ml_ms_count25M(11), ZN => ml_ms_cnt_n_20);
  ml_ms_cnt_count_reg_9 : DFKCNQD1BWP7T port map(CN => ml_ms_cnt_n_23, CP => CTS_288, D => FE_PHN496_ml_ms_cnt_n_17, Q => ml_ms_count25M(9));
  ml_ms_cnt_g230 : MOAI22D0BWP7T port map(A1 => ml_ms_cnt_n_16, A2 => ml_ms_count25M(10), B1 => ml_ms_cnt_n_16, B2 => ml_ms_count25M(10), ZN => ml_ms_cnt_n_19);
  ml_ms_cnt_g231 : IND2D1BWP7T port map(A1 => ml_ms_cnt_n_16, B1 => ml_ms_count25M(10), ZN => ml_ms_cnt_n_18);
  ml_ms_cnt_count_reg_8 : DFKCNQD1BWP7T port map(CN => ml_ms_cnt_n_23, CP => CTS_288, D => FE_PHN495_ml_ms_cnt_n_15, Q => ml_ms_count25M(8));
  ml_ms_cnt_g233 : MOAI22D0BWP7T port map(A1 => ml_ms_cnt_n_14, A2 => ml_ms_count25M(9), B1 => ml_ms_cnt_n_14, B2 => ml_ms_count25M(9), ZN => ml_ms_cnt_n_17);
  ml_ms_cnt_g234 : IND2D1BWP7T port map(A1 => ml_ms_cnt_n_14, B1 => ml_ms_count25M(9), ZN => ml_ms_cnt_n_16);
  ml_ms_cnt_count_reg_7 : DFKCNQD1BWP7T port map(CN => ml_ms_cnt_n_23, CP => CTS_322, D => ml_ms_cnt_n_13, Q => FE_PHN436_ml_ms_count25M_7);
  ml_ms_cnt_g236 : MOAI22D0BWP7T port map(A1 => ml_ms_cnt_n_12, A2 => ml_ms_count25M(8), B1 => ml_ms_cnt_n_12, B2 => ml_ms_count25M(8), ZN => ml_ms_cnt_n_15);
  ml_ms_cnt_g237 : IND2D1BWP7T port map(A1 => ml_ms_cnt_n_12, B1 => ml_ms_count25M(8), ZN => ml_ms_cnt_n_14);
  ml_ms_cnt_count_reg_6 : DFKCNQD1BWP7T port map(CN => ml_ms_cnt_n_11, CP => CTS_322, D => ml_ms_cnt_n_23, Q => ml_ms_count25M(6));
  ml_ms_cnt_g239 : MOAI22D0BWP7T port map(A1 => FE_PHN472_ml_ms_cnt_n_10, A2 => ml_ms_count25M(7), B1 => FE_PHN472_ml_ms_cnt_n_10, B2 => ml_ms_count25M(7), ZN => ml_ms_cnt_n_13);
  ml_ms_cnt_g240 : IND2D1BWP7T port map(A1 => FE_PHN472_ml_ms_cnt_n_10, B1 => ml_ms_count25M(7), ZN => ml_ms_cnt_n_12);
  ml_ms_cnt_count_reg_5 : DFKCNQD1BWP7T port map(CN => FE_PHN507_ml_ms_cnt_n_9, CP => CTS_322, D => ml_ms_cnt_n_23, Q => FE_PHN439_ml_ms_count25M_5);
  ml_ms_cnt_g242 : MOAI22D0BWP7T port map(A1 => ml_ms_cnt_n_8, A2 => FE_PHN415_ml_ms_count25M_6, B1 => ml_ms_cnt_n_8, B2 => FE_PHN415_ml_ms_count25M_6, ZN => FE_PHN474_ml_ms_cnt_n_11);
  ml_ms_cnt_g243 : IND2D1BWP7T port map(A1 => ml_ms_cnt_n_8, B1 => FE_PHN415_ml_ms_count25M_6, ZN => ml_ms_cnt_n_10);
  ml_ms_cnt_count_reg_4 : DFKCNQD1BWP7T port map(CN => FE_PHN508_ml_ms_cnt_n_7, CP => CTS_322, D => ml_ms_cnt_n_23, Q => ml_ms_count25M(4));
  ml_ms_cnt_g245 : MOAI22D0BWP7T port map(A1 => ml_ms_cnt_n_6, A2 => ml_ms_count25M(5), B1 => ml_ms_cnt_n_6, B2 => ml_ms_count25M(5), ZN => ml_ms_cnt_n_9);
  ml_ms_cnt_g246 : IND2D1BWP7T port map(A1 => ml_ms_cnt_n_6, B1 => ml_ms_count25M(5), ZN => ml_ms_cnt_n_8);
  ml_ms_cnt_count_reg_3 : DFKCNQD1BWP7T port map(CN => ml_ms_cnt_n_5, CP => CTS_322, D => ml_ms_cnt_n_23, Q => FE_PHN503_ml_ms_count25M_3);
  ml_ms_cnt_g248 : MOAI22D0BWP7T port map(A1 => ml_ms_cnt_n_4, A2 => FE_PHN437_ml_ms_count25M_4, B1 => ml_ms_cnt_n_4, B2 => FE_PHN437_ml_ms_count25M_4, ZN => ml_ms_cnt_n_7);
  ml_ms_cnt_g249 : IND2D1BWP7T port map(A1 => ml_ms_cnt_n_4, B1 => FE_PHN437_ml_ms_count25M_4, ZN => ml_ms_cnt_n_6);
  ml_ms_cnt_count_reg_2 : DFKCNQD1BWP7T port map(CN => ml_ms_cnt_n_3, CP => CTS_322, D => ml_ms_cnt_n_23, Q => FE_PHN408_ml_ms_count25M_2);
  ml_ms_cnt_g251 : MOAI22D0BWP7T port map(A1 => ml_ms_cnt_n_2, A2 => ml_ms_count25M(3), B1 => ml_ms_cnt_n_2, B2 => ml_ms_count25M(3), ZN => ml_ms_cnt_n_5);
  ml_ms_cnt_g252 : IND2D1BWP7T port map(A1 => ml_ms_cnt_n_2, B1 => ml_ms_count25M(3), ZN => ml_ms_cnt_n_4);
  ml_ms_cnt_count_reg_1 : EDFKCND1BWP7T port map(CN => ml_ms_cnt_n_23, CP => CTS_322, D => FE_PHN447_ml_ms_cnt_count_1, E => ml_ms_cnt_count(0), Q => UNCONNECTED16, QN => ml_ms_cnt_count(1));
  ml_ms_cnt_g254 : MOAI22D0BWP7T port map(A1 => ml_ms_cnt_n_1, A2 => ml_ms_count25M(2), B1 => ml_ms_cnt_n_1, B2 => ml_ms_count25M(2), ZN => ml_ms_cnt_n_3);
  ml_ms_cnt_g255 : IND2D1BWP7T port map(A1 => ml_ms_cnt_n_1, B1 => ml_ms_count25M(2), ZN => ml_ms_cnt_n_2);
  ml_ms_cnt_g257 : IND2D1BWP7T port map(A1 => FE_PHN447_ml_ms_cnt_count_1, B1 => ml_ms_cnt_count(0), ZN => ml_ms_cnt_n_1);
  ml_ms_cnt_count_reg_0 : DFKCND1BWP7T port map(CN => FE_PHN396_ml_ms_cnt_n_0, CP => CTS_322, D => ml_ms_cnt_n_23, Q => FE_PHN378_ml_ms_cnt_count_0, QN => ml_ms_cnt_n_0);
  ml_il_color1_output_color_reg_0 : LHQD1BWP7T port map(D => ml_il_color1_n_18, E => ml_handshake_mouse_out, Q => sig_output_color(0));
  ml_il_color1_output_color_reg_2 : LHQD1BWP7T port map(D => ml_il_color1_n_17, E => ml_handshake_mouse_out, Q => sig_output_color(2));
  ml_il_color1_g273 : IOA21D0BWP7T port map(A1 => ml_il_color1_n_22, A2 => ml_il_color1_state(0), B => ml_il_color1_n_21, ZN => ml_il_color1_n_18);
  ml_il_color1_g274 : OAI21D0BWP7T port map(A1 => ml_il_color1_n_15, A2 => ml_il_color1_state(0), B => ml_il_color1_n_23, ZN => ml_il_color1_n_17);
  ml_il_color1_output_color_reg_1 : LHQD1BWP7T port map(D => ml_il_color1_n_16, E => ml_handshake_mouse_out, Q => sig_output_color(1));
  ml_il_color1_rescount_reg : DFKCNQD1BWP7T port map(CN => ml_il_color1_n_14, CP => CTS_322, D => FE_PHN358_ml_buttons_mouse_3, Q => sig_rescount);
  ml_il_color1_g277 : ND2D0BWP7T port map(A1 => ml_il_color1_n_22, A2 => ml_il_color1_n_21, ZN => ml_il_color1_n_16);
  ml_il_color1_draw_reg : DFQD1BWP7T port map(CP => CTS_288, D => FE_PHN381_ml_buttons_mouse_4, Q => sig_draw);
  ml_il_color1_g280 : IND2D0BWP7T port map(A1 => ml_il_color1_state(1), B1 => ml_il_color1_state(2), ZN => ml_il_color1_n_21);
  ml_il_color1_g281 : INVD0BWP7T port map(I => ml_il_color1_n_15, ZN => ml_il_color1_n_20);
  ml_il_color1_g282 : ND2D0BWP7T port map(A1 => ml_il_color1_state(2), A2 => ml_il_color1_state(1), ZN => ml_il_color1_n_23);
  ml_il_color1_g283 : NR2D0BWP7T port map(A1 => ml_il_color1_state(1), A2 => ml_il_color1_state(2), ZN => ml_il_color1_n_15);
  ml_il_color1_g284 : IND2D0BWP7T port map(A1 => ml_il_color1_state(2), B1 => ml_il_color1_state(1), ZN => ml_il_color1_n_22);
  ml_il_color1_g285 : CKND1BWP7T port map(I => sig_countlow, ZN => ml_il_color1_n_14);
  ml_il_color1_next_state_reg_0 : LHQD1BWP7T port map(D => ml_il_color1_n_12, E => ml_handshake_mouse_out, Q => ml_il_color1_next_state(0));
  ml_il_color1_next_state_reg_1 : LHQD1BWP7T port map(D => ml_il_color1_n_11, E => ml_handshake_mouse_out, Q => ml_il_color1_next_state(1));
  ml_il_color1_g439 : AO22D0BWP7T port map(A1 => ml_il_color1_n_9, A2 => ml_il_color1_state(0), B1 => ml_buttons_mouse(2), B2 => ml_il_color1_n_6, Z => ml_il_color1_n_12);
  ml_il_color1_next_state_reg_2 : LHQD1BWP7T port map(D => ml_il_color1_n_10, E => ml_handshake_mouse_out, Q => ml_il_color1_next_state(2));
  ml_il_color1_g441 : OAI211D0BWP7T port map(A1 => ml_buttons_mouse(2), A2 => ml_il_color1_n_22, B => ml_il_color1_n_8, C => ml_il_color1_n_23, ZN => ml_il_color1_n_11);
  ml_il_color1_g442 : OR3D0BWP7T port map(A1 => ml_il_color1_n_4, A2 => ml_il_color1_n_5, A3 => ml_il_color1_n_7, Z => ml_il_color1_n_10);
  ml_il_color1_g443 : IND3D0BWP7T port map(A1 => ml_il_color1_n_7, B1 => ml_il_color1_n_20, B2 => ml_il_color1_n_22, ZN => ml_il_color1_n_9);
  ml_il_color1_g444 : ND3D0BWP7T port map(A1 => ml_il_color1_n_3, A2 => ml_il_color1_state(0), A3 => ml_buttons_mouse(2), ZN => ml_il_color1_n_8);
  ml_il_color1_state_reg_1 : DFKCNQD1BWP7T port map(CN => ml_il_color1_next_state(1), CP => CTS_288, D => FE_DBTN0_reset, Q => ml_il_color1_state(1));
  ml_il_color1_state_reg_2 : DFKCNQD1BWP7T port map(CN => ml_il_color1_next_state(2), CP => CTS_288, D => FE_DBTN0_reset, Q => ml_il_color1_state(2));
  ml_il_color1_g447 : IND2D0BWP7T port map(A1 => ml_il_color1_n_4, B1 => ml_il_color1_n_20, ZN => ml_il_color1_n_6);
  ml_il_color1_g448 : OAI22D0BWP7T port map(A1 => ml_il_color1_n_21, A2 => ml_il_color1_n_1, B1 => ml_il_color1_n_22, B2 => ml_il_color1_n_0, ZN => ml_il_color1_n_5);
  ml_il_color1_g449 : AOI21D0BWP7T port map(A1 => ml_il_color1_n_21, A2 => ml_il_color1_n_23, B => ml_buttons_mouse(2), ZN => ml_il_color1_n_7);
  ml_il_color1_g450 : NR2D0BWP7T port map(A1 => ml_il_color1_n_23, A2 => ml_il_color1_state(0), ZN => ml_il_color1_n_4);
  ml_il_color1_g451 : ND2D0BWP7T port map(A1 => ml_il_color1_n_21, A2 => ml_il_color1_n_20, ZN => ml_il_color1_n_3);
  ml_il_color1_g454 : INVD0BWP7T port map(I => ml_buttons_mouse(2), ZN => ml_il_color1_n_0);
  ml_il_color1_state_reg_0 : DFKCND1BWP7T port map(CN => ml_il_color1_next_state(0), CP => CTS_288, D => FE_DBTN0_reset, Q => ml_il_color1_state(0), QN => ml_il_color1_n_1);
  gl_vgd_g1603 : OR2D1BWP7T port map(A1 => gl_vgd_n_83, A2 => gl_vgd_horizontal(8), Z => FE_OFN34_H);
  gl_vgd_g1604 : IND4D0BWP7T port map(A1 => gl_vgd_n_79, B1 => gl_vgd_horizontal(7), B2 => gl_vgd_horizontal(9), B3 => gl_vgd_n_81, ZN => gl_vgd_n_83);
  gl_vgd_g1605 : NR4D0BWP7T port map(A1 => gl_vgd_n_78, A2 => gl_vgd_n_74, A3 => gl_vgd_horizontal(4), A4 => gl_vgd_horizontal(1), ZN => gl_sig_scale_h);
  gl_vgd_g1606 : CKAN2D8BWP7T port map(A1 => gl_vgd_n_82, A2 => gl_sig_red, Z => R);
  gl_vgd_g1607 : ND2D5BWP7T port map(A1 => gl_vgd_n_82, A2 => gl_vgd_n_67, ZN => G);
  gl_vgd_g1608 : CKAN2D8BWP7T port map(A1 => gl_vgd_n_82, A2 => gl_sig_blue, Z => B);
  gl_vgd_g1609 : OR3XD1BWP7T port map(A1 => gl_vgd_vertical(9), A2 => gl_vgd_n_73, A3 => gl_vgd_n_80, Z => FE_OFN35_V);
  gl_vgd_g1610 : IINR4D0BWP7T port map(A1 => gl_vgd_n_77, A2 => gl_vgd_n_73, B1 => gl_vgd_vertical(1), B2 => gl_vgd_vertical(9), ZN => gl_sig_scale_v);
  gl_vgd_g1611 : INR3D0BWP7T port map(A1 => gl_vgd_n_73, B1 => gl_vgd_vertical(9), B2 => gl_vgd_n_78, ZN => gl_vgd_n_82);
  gl_vgd_g1612 : OAI211D1BWP7T port map(A1 => gl_vgd_n_72, A2 => gl_vgd_n_75, B => gl_vgd_horizontal(6), C => gl_vgd_horizontal(5), ZN => gl_vgd_n_81);
  gl_vgd_g1613 : IND4D0BWP7T port map(A1 => gl_vgd_vertical(4), B1 => gl_vgd_vertical(3), B2 => gl_vgd_n_69, B3 => gl_vgd_n_71, ZN => gl_vgd_n_80);
  gl_vgd_g1614 : AOI211XD0BWP7T port map(A1 => gl_vgd_n_75, A2 => gl_vgd_n_68, B => gl_vgd_horizontal(6), C => gl_vgd_horizontal(5), ZN => gl_vgd_n_79);
  gl_vgd_g1615 : IND2D1BWP7T port map(A1 => gl_vgd_horizontal(9), B1 => gl_vgd_n_76, ZN => gl_vgd_n_78);
  gl_vgd_g1616 : NR3D0BWP7T port map(A1 => gl_vgd_n_69, A2 => gl_vgd_vertical(4), A3 => gl_vgd_vertical(3), ZN => gl_vgd_n_77);
  gl_vgd_g1617 : ND4D0BWP7T port map(A1 => gl_vgd_horizontal(5), A2 => gl_vgd_horizontal(6), A3 => gl_vgd_horizontal(7), A4 => gl_vgd_horizontal(8), ZN => gl_vgd_n_76);
  gl_vgd_g1618 : IND2D1BWP7T port map(A1 => gl_vgd_horizontal(0), B1 => gl_vgd_n_70, ZN => gl_vgd_n_74);
  gl_vgd_g1619 : INR2D1BWP7T port map(A1 => gl_vgd_horizontal(4), B1 => gl_vgd_n_70, ZN => gl_vgd_n_75);
  gl_vgd_g1620 : AN3D1BWP7T port map(A1 => gl_vgd_horizontal(4), A2 => gl_vgd_horizontal(1), A3 => gl_vgd_horizontal(0), Z => gl_vgd_n_72);
  gl_vgd_g1621 : MUX2ND0BWP7T port map(I0 => gl_vgd_vertical(0), I1 => gl_vgd_vertical(2), S => gl_vgd_vertical(1), ZN => gl_vgd_n_71);
  gl_vgd_g1622 : ND4D0BWP7T port map(A1 => gl_vgd_vertical(5), A2 => gl_vgd_vertical(6), A3 => gl_vgd_vertical(8), A4 => gl_vgd_vertical(7), ZN => gl_vgd_n_73);
  gl_vgd_g1623 : NR2XD0BWP7T port map(A1 => gl_vgd_horizontal(3), A2 => gl_vgd_horizontal(2), ZN => gl_vgd_n_70);
  gl_vgd_g1624 : OR2D1BWP7T port map(A1 => gl_vgd_horizontal(3), A2 => gl_vgd_horizontal(1), Z => gl_vgd_n_68);
  gl_vgd_g1625 : OR2D1BWP7T port map(A1 => gl_vgd_vertical(2), A2 => gl_vgd_vertical(0), Z => gl_vgd_n_69);
  gl_vgd_scale_horizontal_reg_2 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_288, D => FE_PHN448_gl_vgd_horizontal_counter_2, Q => gl_vgd_horizontal(2));
  gl_vgd_vertical_reg_3 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_288, D => FE_PHN419_gl_vgd_vertical_counter_3, Q => gl_vgd_vertical(3));
  gl_vgd_scale_horizontal_reg_3 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_288, D => FE_PHN445_gl_vgd_horizontal_counter_3, Q => gl_vgd_horizontal(3));
  gl_vgd_vertical_reg_0 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_288, D => FE_PHN412_gl_vgd_vertical_counter_0, Q => gl_vgd_vertical(0));
  gl_vgd_vertical_reg_2 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_288, D => FE_PHN409_gl_vgd_vertical_counter_2, Q => gl_vgd_vertical(2));
  gl_vgd_horizontal_reg_7 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_288, D => gl_vgd_horizontal_counter(7), Q => gl_vgd_horizontal(7));
  gl_vgd_vertical_reg_4 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_288, D => gl_vgd_vertical_counter(4), Q => gl_vgd_vertical(4));
  gl_vgd_scale_horizontal_reg_4 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_288, D => FE_PHN449_gl_vgd_horizontal_counter_4, Q => gl_vgd_horizontal(4));
  gl_vgd_horizontal_reg_5 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_288, D => FE_PHN446_gl_vgd_horizontal_counter_5, Q => gl_vgd_horizontal(5));
  gl_vgd_scale_horizontal_reg_6 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_288, D => FE_PHN450_gl_vgd_horizontal_counter_6, Q => gl_vgd_horizontal(6));
  gl_vgd_vertical_reg_5 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_288, D => gl_vgd_vertical_counter(5), Q => gl_vgd_vertical(5));
  gl_vgd_scale_vertical_reg_6 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_288, D => gl_vgd_vertical_counter(6), Q => gl_vgd_vertical(6));
  gl_vgd_scale_vertical_reg_8 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_288, D => gl_vgd_vertical_counter(8), Q => gl_vgd_vertical(8));
  gl_vgd_scale_vertical_reg_7 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_288, D => gl_vgd_vertical_counter(7), Q => gl_vgd_vertical(7));
  gl_vgd_horizontal_reg_9 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_288, D => gl_vgd_horizontal_counter(9), Q => gl_vgd_horizontal(9));
  gl_vgd_scale_horizontal_reg_8 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_288, D => FE_PHN451_gl_vgd_horizontal_counter_8, Q => gl_vgd_horizontal(8));
  gl_vgd_horizontal_reg_0 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_288, D => gl_vgd_horizontal_counter(0), Q => gl_vgd_horizontal(0));
  gl_vgd_vertical_reg_1 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_288, D => gl_vgd_vertical_counter(1), Q => gl_vgd_vertical(1));
  gl_vgd_scale_horizontal_reg_1 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_288, D => gl_vgd_horizontal_counter(1), Q => gl_vgd_horizontal(1));
  gl_vgd_scale_vertical_reg_9 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_288, D => gl_vgd_vertical_counter(9), Q => gl_vgd_vertical(9));
  gl_vgd_g1646 : INVD1BWP7T port map(I => gl_sig_green, ZN => gl_vgd_n_67);
  gl_vgd_horizontal_counter_reg_0 : DFKCNQD1BWP7T port map(CN => gl_vgd_n_6, CP => CTS_288, D => gl_vgd_n_41, Q => FE_PHN435_gl_vgd_horizontal_counter_0);
  gl_vgd_horizontal_counter_reg_1 : DFKCNQD1BWP7T port map(CN => gl_vgd_n_19, CP => CTS_288, D => gl_vgd_n_41, Q => FE_PHN444_gl_vgd_horizontal_counter_1);
  gl_vgd_horizontal_counter_reg_2 : DFKCNQD1BWP7T port map(CN => gl_vgd_n_24, CP => CTS_288, D => gl_vgd_n_41, Q => gl_vgd_horizontal_counter(2));
  gl_vgd_horizontal_counter_reg_3 : DFKCNQD1BWP7T port map(CN => gl_vgd_n_29, CP => CTS_288, D => gl_vgd_n_41, Q => gl_vgd_horizontal_counter(3));
  gl_vgd_horizontal_counter_reg_4 : DFKCNQD1BWP7T port map(CN => gl_vgd_n_32, CP => CTS_288, D => gl_vgd_n_41, Q => gl_vgd_horizontal_counter(4));
  gl_vgd_horizontal_counter_reg_5 : DFKCNQD1BWP7T port map(CN => gl_vgd_n_37, CP => CTS_288, D => gl_vgd_n_41, Q => gl_vgd_horizontal_counter(5));
  gl_vgd_horizontal_counter_reg_6 : DFKCNQD1BWP7T port map(CN => gl_vgd_n_46, CP => CTS_288, D => gl_vgd_n_41, Q => gl_vgd_horizontal_counter(6));
  gl_vgd_horizontal_counter_reg_7 : DFKCNQD1BWP7T port map(CN => gl_vgd_n_56, CP => CTS_288, D => gl_vgd_n_41, Q => FE_PHN453_gl_vgd_horizontal_counter_7);
  gl_vgd_horizontal_counter_reg_8 : DFKCNQD1BWP7T port map(CN => gl_vgd_n_41, CP => CTS_288, D => gl_vgd_n_62, Q => gl_vgd_horizontal_counter(8));
  gl_vgd_horizontal_counter_reg_9 : DFKCNQD1BWP7T port map(CN => gl_vgd_n_41, CP => CTS_288, D => gl_vgd_n_65, Q => FE_PHN432_gl_vgd_horizontal_counter_9);
  gl_vgd_vertical_counter_reg_0 : DFXQD1BWP7T port map(CP => CTS_288, DA => gl_vgd_n_44, DB => gl_vgd_n_43, Q => gl_vgd_vertical_counter(0), SA => FE_PHN412_gl_vgd_vertical_counter_0);
  gl_vgd_vertical_counter_reg_1 : DFQD1BWP7T port map(CP => CTS_288, D => gl_vgd_n_51, Q => FE_PHN410_gl_vgd_vertical_counter_1);
  gl_vgd_vertical_counter_reg_2 : DFQD1BWP7T port map(CP => CTS_288, D => gl_vgd_n_52, Q => gl_vgd_vertical_counter(2));
  gl_vgd_vertical_counter_reg_3 : DFQD1BWP7T port map(CP => CTS_288, D => gl_vgd_n_49, Q => gl_vgd_vertical_counter(3));
  gl_vgd_vertical_counter_reg_4 : DFQD1BWP7T port map(CP => CTS_288, D => gl_vgd_n_54, Q => FE_PHN418_gl_vgd_vertical_counter_4);
  gl_vgd_vertical_counter_reg_5 : DFQD1BWP7T port map(CP => CTS_288, D => gl_vgd_n_53, Q => FE_PHN423_gl_vgd_vertical_counter_5);
  gl_vgd_vertical_counter_reg_6 : DFQD1BWP7T port map(CP => CTS_288, D => gl_vgd_n_50, Q => FE_PHN421_gl_vgd_vertical_counter_6);
  gl_vgd_vertical_counter_reg_7 : DFQD1BWP7T port map(CP => CTS_288, D => gl_vgd_n_57, Q => FE_PHN433_gl_vgd_vertical_counter_7);
  gl_vgd_vertical_counter_reg_9 : DFQD1BWP7T port map(CP => CTS_288, D => FE_PHN468_gl_vgd_n_64, Q => FE_PHN442_gl_vgd_vertical_counter_9);
  gl_vgd_g1735 : MOAI22D0BWP7T port map(A1 => gl_vgd_n_63, A2 => gl_vgd_n_14, B1 => gl_vgd_n_63, B2 => gl_vgd_n_14, ZN => gl_vgd_n_65);
  gl_vgd_g1738 : AO22D0BWP7T port map(A1 => gl_vgd_n_58, A2 => gl_vgd_vertical_counter(9), B1 => gl_vgd_n_60, B2 => gl_vgd_n_43, Z => gl_vgd_n_64);
  gl_vgd_g1739 : HA1D0BWP7T port map(A => gl_vgd_n_11, B => gl_vgd_n_55, CO => gl_vgd_n_63, S => gl_vgd_n_62);
  gl_vgd_g1740 : AO21D0BWP7T port map(A1 => gl_vgd_n_58, A2 => gl_vgd_vertical_counter(8), B => gl_vgd_n_59, Z => gl_vgd_n_61);
  gl_vgd_g1742 : OAI31D0BWP7T port map(A1 => gl_vgd_vertical_counter(9), A2 => gl_vgd_n_2, A3 => gl_vgd_n_47, B => gl_vgd_n_15, ZN => gl_vgd_n_60);
  gl_vgd_g1744 : NR3D0BWP7T port map(A1 => gl_vgd_n_42, A2 => gl_vgd_n_47, A3 => gl_vgd_vertical_counter(8), ZN => gl_vgd_n_59);
  gl_vgd_g1745 : MOAI22D0BWP7T port map(A1 => gl_vgd_n_42, A2 => gl_vgd_n_48, B1 => gl_vgd_n_44, B2 => gl_vgd_vertical_counter(7), ZN => gl_vgd_n_57);
  gl_vgd_g1746 : AO21D0BWP7T port map(A1 => gl_vgd_n_43, A2 => gl_vgd_n_47, B => gl_vgd_n_44, Z => gl_vgd_n_58);
  gl_vgd_g1747 : HA1D0BWP7T port map(A => gl_vgd_n_13, B => gl_vgd_n_45, CO => gl_vgd_n_55, S => gl_vgd_n_56);
  gl_vgd_g1755 : MOAI22D0BWP7T port map(A1 => gl_vgd_n_42, A2 => gl_vgd_n_30, B1 => gl_vgd_n_44, B2 => gl_vgd_vertical_counter(4), ZN => gl_vgd_n_54);
  gl_vgd_g1756 : MOAI22D0BWP7T port map(A1 => gl_vgd_n_42, A2 => gl_vgd_n_34, B1 => gl_vgd_n_44, B2 => gl_vgd_vertical_counter(5), ZN => gl_vgd_n_53);
  gl_vgd_g1758 : MOAI22D0BWP7T port map(A1 => gl_vgd_n_42, A2 => gl_vgd_n_20, B1 => gl_vgd_n_44, B2 => FE_PHN409_gl_vgd_vertical_counter_2, ZN => gl_vgd_n_52);
  gl_vgd_g1759 : MOAI22D0BWP7T port map(A1 => gl_vgd_n_42, A2 => gl_vgd_n_0, B1 => gl_vgd_n_44, B2 => gl_vgd_vertical_counter(1), ZN => gl_vgd_n_51);
  gl_vgd_g1760 : MOAI22D0BWP7T port map(A1 => gl_vgd_n_42, A2 => gl_vgd_n_39, B1 => gl_vgd_n_44, B2 => gl_vgd_vertical_counter(6), ZN => gl_vgd_n_50);
  gl_vgd_g1761 : MOAI22D0BWP7T port map(A1 => gl_vgd_n_42, A2 => gl_vgd_n_25, B1 => gl_vgd_n_44, B2 => FE_PHN419_gl_vgd_vertical_counter_3, ZN => gl_vgd_n_49);
  gl_vgd_g1765 : MAOI22D0BWP7T port map(A1 => gl_vgd_n_38, A2 => gl_vgd_vertical_counter(7), B1 => gl_vgd_n_38, B2 => gl_vgd_vertical_counter(7), ZN => gl_vgd_n_48);
  gl_vgd_g1769 : HA1D0BWP7T port map(A => gl_vgd_n_12, B => gl_vgd_n_36, CO => gl_vgd_n_45, S => gl_vgd_n_46);
  gl_vgd_g1770 : IND2D1BWP7T port map(A1 => gl_vgd_n_38, B1 => gl_vgd_vertical_counter(7), ZN => gl_vgd_n_47);
  gl_vgd_g1771 : INVD1BWP7T port map(I => gl_vgd_n_43, ZN => gl_vgd_n_42);
  gl_vgd_g1772 : NR2D1BWP7T port map(A1 => gl_vgd_n_40, A2 => FE_OFN31_reset, ZN => gl_vgd_n_44);
  gl_vgd_g1773 : NR2XD0BWP7T port map(A1 => gl_vgd_n_41, A2 => gl_vgd_n_26, ZN => gl_vgd_n_43);
  gl_vgd_g1774 : INVD1BWP7T port map(I => gl_vgd_n_41, ZN => gl_vgd_n_40);
  gl_vgd_g1775 : IND3D1BWP7T port map(A1 => gl_vgd_n_13, B1 => gl_vgd_n_11, B2 => gl_vgd_n_35, ZN => gl_vgd_n_41);
  gl_vgd_g1776 : MAOI22D0BWP7T port map(A1 => gl_vgd_n_31, A2 => gl_vgd_vertical_counter(6), B1 => gl_vgd_n_31, B2 => gl_vgd_vertical_counter(6), ZN => gl_vgd_n_39);
  gl_vgd_g1777 : HA1D0BWP7T port map(A => gl_vgd_n_8, B => gl_vgd_n_33, CO => gl_vgd_n_36, S => gl_vgd_n_37);
  gl_vgd_g1778 : IND2D1BWP7T port map(A1 => gl_vgd_n_31, B1 => gl_vgd_vertical_counter(6), ZN => gl_vgd_n_38);
  gl_vgd_g1779 : INR4D0BWP7T port map(A1 => gl_vgd_n_33, B1 => gl_vgd_n_14, B2 => gl_vgd_n_8, B3 => gl_vgd_n_12, ZN => gl_vgd_n_35);
  gl_vgd_g1780 : MAOI22D0BWP7T port map(A1 => gl_vgd_n_27, A2 => gl_vgd_vertical_counter(5), B1 => gl_vgd_n_27, B2 => gl_vgd_vertical_counter(5), ZN => gl_vgd_n_34);
  gl_vgd_g1781 : HA1D0BWP7T port map(A => gl_vgd_n_10, B => gl_vgd_n_28, CO => gl_vgd_n_33, S => gl_vgd_n_32);
  gl_vgd_g1782 : IND2D1BWP7T port map(A1 => gl_vgd_n_27, B1 => gl_vgd_vertical_counter(5), ZN => gl_vgd_n_31);
  gl_vgd_g1783 : MAOI22D0BWP7T port map(A1 => gl_vgd_n_22, A2 => gl_vgd_vertical_counter(4), B1 => gl_vgd_n_22, B2 => gl_vgd_vertical_counter(4), ZN => gl_vgd_n_30);
  gl_vgd_g1784 : HA1D0BWP7T port map(A => gl_vgd_n_4, B => gl_vgd_n_23, CO => gl_vgd_n_28, S => gl_vgd_n_29);
  gl_vgd_g1785 : IND2D1BWP7T port map(A1 => gl_vgd_n_22, B1 => gl_vgd_vertical_counter(4), ZN => gl_vgd_n_27);
  gl_vgd_g1786 : NR4D0BWP7T port map(A1 => gl_vgd_n_21, A2 => gl_vgd_vertical_counter(7), A3 => gl_vgd_vertical_counter(6), A4 => gl_vgd_vertical_counter(5), ZN => gl_vgd_n_26);
  gl_vgd_g1787 : MAOI22D0BWP7T port map(A1 => gl_vgd_n_17, A2 => FE_PHN419_gl_vgd_vertical_counter_3, B1 => gl_vgd_n_17, B2 => FE_PHN419_gl_vgd_vertical_counter_3, ZN => gl_vgd_n_25);
  gl_vgd_g1788 : HA1D0BWP7T port map(A => gl_vgd_n_3, B => gl_vgd_n_18, CO => gl_vgd_n_23, S => gl_vgd_n_24);
  gl_vgd_g1789 : IND2D1BWP7T port map(A1 => gl_vgd_n_17, B1 => FE_PHN419_gl_vgd_vertical_counter_3, ZN => gl_vgd_n_22);
  gl_vgd_g1790 : IND4D0BWP7T port map(A1 => gl_vgd_vertical_counter(4), B1 => FE_PHN409_gl_vgd_vertical_counter_2, B2 => FE_PHN419_gl_vgd_vertical_counter_3, B3 => gl_vgd_n_16, ZN => gl_vgd_n_21);
  gl_vgd_g1791 : MAOI22D0BWP7T port map(A1 => gl_vgd_n_9, A2 => FE_PHN409_gl_vgd_vertical_counter_2, B1 => gl_vgd_n_9, B2 => FE_PHN409_gl_vgd_vertical_counter_2, ZN => gl_vgd_n_20);
  gl_vgd_g1792 : HA1D0BWP7T port map(A => gl_vgd_n_7, B => gl_vgd_n_5, CO => gl_vgd_n_18, S => gl_vgd_n_19);
  gl_vgd_g1793 : IND2D1BWP7T port map(A1 => gl_vgd_n_9, B1 => FE_PHN409_gl_vgd_vertical_counter_2, ZN => gl_vgd_n_17);
  gl_vgd_g1794 : NR3D0BWP7T port map(A1 => gl_vgd_n_15, A2 => gl_vgd_vertical_counter(1), A3 => FE_PHN412_gl_vgd_vertical_counter_0, ZN => gl_vgd_n_16);
  gl_vgd_g1796 : ND2D1BWP7T port map(A1 => gl_vgd_n_2, A2 => gl_vgd_vertical_counter(9), ZN => gl_vgd_n_15);
  gl_vgd_g1797 : ND2D1BWP7T port map(A1 => gl_vgd_horizontal_counter(9), A2 => FE_DBTN0_reset, ZN => gl_vgd_n_14);
  gl_vgd_g1798 : INR2XD0BWP7T port map(A1 => FE_PHN449_gl_vgd_horizontal_counter_4, B1 => FE_OFN31_reset, ZN => gl_vgd_n_10);
  gl_vgd_g1799 : INR2D1BWP7T port map(A1 => gl_vgd_horizontal_counter(7), B1 => FE_OFN31_reset, ZN => gl_vgd_n_13);
  gl_vgd_g1800 : INR2D1BWP7T port map(A1 => FE_PHN450_gl_vgd_horizontal_counter_6, B1 => FE_OFN31_reset, ZN => gl_vgd_n_12);
  gl_vgd_g1801 : INR2D1BWP7T port map(A1 => FE_PHN451_gl_vgd_horizontal_counter_8, B1 => FE_OFN31_reset, ZN => gl_vgd_n_11);
  gl_vgd_g1802 : INVD0BWP7T port map(I => gl_vgd_n_6, ZN => gl_vgd_n_7);
  gl_vgd_g1803 : CKAN2D1BWP7T port map(A1 => gl_vgd_horizontal_counter(1), A2 => FE_DBTN0_reset, Z => gl_vgd_n_5);
  gl_vgd_g1804 : ND2D1BWP7T port map(A1 => gl_vgd_vertical_counter(1), A2 => FE_PHN412_gl_vgd_vertical_counter_0, ZN => gl_vgd_n_9);
  gl_vgd_g1805 : CKAN2D1BWP7T port map(A1 => FE_PHN445_gl_vgd_horizontal_counter_3, A2 => FE_DBTN0_reset, Z => gl_vgd_n_4);
  gl_vgd_g1806 : CKAN2D1BWP7T port map(A1 => FE_PHN448_gl_vgd_horizontal_counter_2, A2 => FE_DBTN0_reset, Z => gl_vgd_n_3);
  gl_vgd_g1807 : AN2D1BWP7T port map(A1 => FE_PHN446_gl_vgd_horizontal_counter_5, A2 => FE_DBTN0_reset, Z => gl_vgd_n_8);
  gl_vgd_g1808 : ND2D1BWP7T port map(A1 => gl_vgd_horizontal_counter(0), A2 => FE_DBTN0_reset, ZN => gl_vgd_n_6);
  gl_vgd_g2 : XNR2D1BWP7T port map(A1 => gl_vgd_vertical_counter(1), A2 => FE_PHN412_gl_vgd_vertical_counter_0, ZN => gl_vgd_n_0);
  gl_vgd_vertical_counter_reg_8 : DFD1BWP7T port map(CP => CTS_288, D => gl_vgd_n_61, Q => FE_PHN359_gl_vgd_vertical_counter_8, QN => gl_vgd_n_2);
  ml_il_x1_g531 : OAI222D0BWP7T port map(A1 => ml_il_x1_n_27, A2 => ml_il_x1_n_6, B1 => ml_il_x1_n_3, B2 => ml_il_x1_cmbsop_sel(1), C1 => ml_il_x1_n_8, C2 => ml_il_x1_n_29, ZN => ml_il_x1_input_register(3));
  ml_il_x1_g532 : MAOI22D0BWP7T port map(A1 => ml_il_x1_n_28, A2 => ml_il_x1_input_register(3), B1 => ml_il_x1_n_28, B2 => ml_il_x1_input_register(3), ZN => ml_il_x1_n_29);
  ml_il_x1_g533 : AO21D0BWP7T port map(A1 => ml_il_x1_n_25, A2 => ml_il_x1_n_17, B => ml_il_x1_n_20, Z => ml_il_x1_n_28);
  ml_il_x1_g534 : MAOI22D0BWP7T port map(A1 => ml_il_x1_n_26, A2 => ml_il_x1_input_register(3), B1 => ml_il_x1_n_26, B2 => ml_il_x1_input_register(3), ZN => ml_il_x1_n_27);
  ml_il_x1_g535 : MOAI22D0BWP7T port map(A1 => ml_il_x1_n_25, A2 => ml_il_x1_n_23, B1 => ml_il_x1_n_25, B2 => ml_il_x1_n_23, ZN => ml_il_x1_n_40);
  ml_il_x1_g536 : MAOI222D1BWP7T port map(A => ml_il_x1_n_24, B => ml_il_x1_n_49, C => ml_mouseX(2), ZN => ml_il_x1_n_26);
  ml_il_x1_g537 : AO21D0BWP7T port map(A1 => ml_il_x1_n_16, A2 => ml_il_x1_n_21, B => ml_il_x1_n_18, Z => ml_il_x1_n_25);
  ml_il_x1_g538 : CKXOR2D0BWP7T port map(A1 => ml_il_x1_n_24, A2 => ml_il_x1_n_23, Z => ml_il_x1_n_39);
  ml_il_x1_g539 : MOAI22D0BWP7T port map(A1 => ml_il_x1_n_22, A2 => ml_il_x1_n_16, B1 => ml_il_x1_n_22, B2 => ml_il_x1_n_16, ZN => ml_il_x1_n_42);
  ml_il_x1_g540 : MOAI22D0BWP7T port map(A1 => ml_il_x1_n_22, A2 => ml_il_x1_n_19, B1 => ml_il_x1_n_22, B2 => ml_il_x1_n_19, ZN => ml_il_x1_n_41);
  ml_il_x1_g541 : MAOI222D1BWP7T port map(A => ml_il_x1_n_19, B => ml_il_x1_n_14, C => ml_il_x1_n_4, ZN => ml_il_x1_n_24);
  ml_il_x1_g542 : IND2D0BWP7T port map(A1 => ml_il_x1_n_20, B1 => ml_il_x1_n_17, ZN => ml_il_x1_n_23);
  ml_il_x1_g543 : OAI21D0BWP7T port map(A1 => ml_il_x1_n_15, A2 => ml_mouseX(0), B => ml_il_x1_n_16, ZN => ml_il_x1_n_43);
  ml_il_x1_g544 : IND2D0BWP7T port map(A1 => ml_il_x1_n_18, B1 => ml_il_x1_n_21, ZN => ml_il_x1_n_22);
  ml_il_x1_g545 : ND2D1BWP7T port map(A1 => ml_il_x1_n_14, A2 => ml_mouseX(1), ZN => ml_il_x1_n_21);
  ml_il_x1_g546 : NR2D0BWP7T port map(A1 => ml_il_x1_n_13, A2 => ml_mouseX(2), ZN => ml_il_x1_n_20);
  ml_il_x1_g547 : ND2D1BWP7T port map(A1 => ml_il_x1_n_47, A2 => ml_mouseX(0), ZN => ml_il_x1_n_19);
  ml_il_x1_g548 : NR2D0BWP7T port map(A1 => ml_il_x1_n_14, A2 => ml_mouseX(1), ZN => ml_il_x1_n_18);
  ml_il_x1_g549 : ND2D1BWP7T port map(A1 => ml_il_x1_n_13, A2 => ml_mouseX(2), ZN => ml_il_x1_n_17);
  ml_il_x1_g550 : ND2D1BWP7T port map(A1 => ml_il_x1_n_15, A2 => ml_mouseX(0), ZN => ml_il_x1_n_16);
  ml_il_x1_g551 : CKND1BWP7T port map(I => ml_il_x1_n_47, ZN => ml_il_x1_n_15);
  ml_il_x1_g553 : INVD1BWP7T port map(I => ml_il_x1_n_48, ZN => ml_il_x1_n_14);
  ml_il_x1_g554 : CKND1BWP7T port map(I => ml_il_x1_n_49, ZN => ml_il_x1_n_13);
  ml_il_x1_g560 : INVD1BWP7T port map(I => ml_il_x1_n_8, ZN => ml_il_x1_n_9);
  ml_il_x1_g561 : ND2D1BWP7T port map(A1 => ml_il_x1_cmbsop_sel(1), A2 => ml_buttons_mouse(0), ZN => ml_il_x1_n_8);
  ml_il_x1_g562 : INVD0BWP7T port map(I => ml_il_x1_n_7, ZN => ml_il_x1_n_6);
  ml_il_x1_g563 : NR2XD0BWP7T port map(A1 => ml_il_x1_n_5, A2 => ml_buttons_mouse(0), ZN => ml_il_x1_n_7);
  ml_il_x1_g564 : INVD1BWP7T port map(I => ml_il_x1_cmbsop_sel(1), ZN => ml_il_x1_n_5);
  ml_il_x1_g565 : INR2D1BWP7T port map(A1 => FE_PHN441_ml_il_x1_state_0, B1 => ml_il_x1_state(1), ZN => ml_il_x1_cmbsop_sel(1));
  ml_il_x1_g566 : INVD0BWP7T port map(I => ml_mouseX(1), ZN => ml_il_x1_n_4);
  ml_il_x1_state_reg_0 : DFQD1BWP7T port map(CP => CTS_322, D => ml_il_x1_n_2, Q => ml_il_x1_state(0));
  ml_il_x1_state_reg_1 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_322, D => ml_il_x1_n_1, Q => FE_PHN431_ml_il_x1_state_1);
  ml_il_x1_g255 : INR4D0BWP7T port map(A1 => ml_handshake_mouse_out, B1 => FE_OFN31_reset, B2 => ml_il_x1_state(1), B3 => FE_PHN441_ml_il_x1_state_0, ZN => ml_il_x1_n_2);
  ml_il_x1_tempx_reg_0 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_322, D => FE_PHN484_ml_il_x1_n_47, Q => FE_PHN513_sig_logic_x_0);
  ml_il_x1_tempx_reg_1 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_322, D => FE_PHN481_ml_il_x1_n_48, Q => FE_PHN512_sig_logic_x_1);
  ml_il_x1_tempx_reg_2 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_322, D => ml_il_x1_n_49, Q => FE_PHN514_sig_logic_x_2);
  ml_il_x1_g260 : AO21D0BWP7T port map(A1 => ml_handshake_mouse_out, A2 => ml_il_x1_state(1), B => ml_il_x1_cmbsop_sel(1), Z => ml_il_x1_n_1);
  ml_il_x1_tempx_reg_3 : DFKCND1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_322, D => FE_PHN497_ml_il_x1_input_register_3, Q => sig_logic_x(3), QN => ml_il_x1_n_3);
  ml_il_x1_g2 : AO222D0BWP7T port map(A1 => ml_il_x1_n_7, A2 => ml_il_x1_n_43, B1 => ml_il_x1_n_9, B2 => ml_il_x1_n_43, C1 => ml_il_x1_n_5, C2 => FE_PHN505_sig_logic_x_0, Z => ml_il_x1_n_47);
  ml_il_x1_g570 : AO222D0BWP7T port map(A1 => ml_il_x1_n_7, A2 => ml_il_x1_n_41, B1 => ml_il_x1_n_9, B2 => ml_il_x1_n_42, C1 => ml_il_x1_n_5, C2 => sig_logic_x(1), Z => ml_il_x1_n_48);
  ml_il_x1_g571 : AO222D0BWP7T port map(A1 => ml_il_x1_n_7, A2 => ml_il_x1_n_39, B1 => ml_il_x1_n_9, B2 => ml_il_x1_n_40, C1 => ml_il_x1_n_5, C2 => sig_logic_x(2), Z => ml_il_x1_n_49);
  ml_ms_mx2_g23 : MUX2D1BWP7T port map(I0 => ml_ms_cntReset25M_main, I1 => ml_ms_cntReset25M_send, S => ml_ms_mux_select_main, Z => ml_ms_cntReset25M);
  ml_ms_ed_reg2_reg : DFQD1BWP7T port map(CP => CTS_322, D => ml_ms_ed_reg1, Q => ml_ms_ed_reg2);
  ml_ms_ed_g224 : NR2XD0BWP7T port map(A1 => ml_ms_ed_n_9, A2 => ml_ms_ed_state(0), ZN => ml_ms_output_edgedet);
  ml_ms_ed_g399 : OAI32D1BWP7T port map(A1 => FE_OFN31_reset, A2 => ml_ms_ed_state(1), A3 => ml_ms_ed_n_5, B1 => ml_ms_ed_n_9, B2 => ml_ms_ed_n_6, ZN => ml_ms_ed_n_8);
  ml_ms_ed_g400 : INVD0BWP7T port map(I => ml_ms_ed_n_6, ZN => ml_ms_ed_n_7);
  ml_ms_ed_g401 : IND2D1BWP7T port map(A1 => FE_OFN31_reset, B1 => ml_ms_ed_n_5, ZN => ml_ms_ed_n_6);
  ml_ms_ed_g402 : OAI31D0BWP7T port map(A1 => FE_PHN361_ml_ms_count_debounce_9, A2 => FE_PHN360_ml_ms_count_debounce_8, A3 => ml_ms_ed_n_4, B => ml_ms_ed_state(0), ZN => FE_PHN456_ml_ms_ed_n_5);
  ml_ms_ed_g403 : OR4D1BWP7T port map(A1 => ml_ms_count_debounce(11), A2 => ml_ms_count_debounce(10), A3 => ml_ms_count_debounce(12), A4 => ml_ms_ed_n_3, Z => ml_ms_ed_n_4);
  ml_ms_ed_g404 : OA31D1BWP7T port map(A1 => FE_PHN377_ml_ms_count_debounce_3, A2 => ml_ms_count_debounce(5), A3 => FE_PHN375_ml_ms_count_debounce_4, B => ml_ms_ed_n_1, Z => ml_ms_ed_n_3);
  ml_ms_ed_g405 : AO211D0BWP7T port map(A1 => ml_ms_ed_n_0, A2 => ml_ms_ed_reg2, B => ml_ms_ed_state(1), C => ml_ms_ed_state(0), Z => ml_ms_ed_n_2);
  ml_ms_ed_g406 : AN2D0BWP7T port map(A1 => ml_ms_count_debounce(6), A2 => ml_ms_count_debounce(7), Z => ml_ms_ed_n_1);
  ml_ms_ed_state_reg_0 : DFKCND1BWP7T port map(CN => FE_PHN467_ml_ms_ed_n_2, CP => CTS_322, D => ml_ms_ed_n_7, Q => ml_ms_ed_state(0), QN => ml_ms_count_debounce_reset);
  ml_ms_ed_state_reg_1 : DFD1BWP7T port map(CP => CTS_322, D => FE_PHN488_ml_ms_ed_n_8, Q => FE_PHN362_ml_ms_ed_state_1, QN => ml_ms_ed_n_9);
  ml_ms_ed_reg1_reg : DFD1BWP7T port map(CP => CTS_322, D => FE_PHN438_clk15k_in, Q => FE_PHN370_ml_ms_ed_reg1, QN => ml_ms_ed_n_0);
  ml_ms_cntD_g71 : INVD1BWP7T port map(I => ml_ms_count_debounce_reset, ZN => ml_ms_cntD_n_23);
  ml_ms_cntD_count_reg_12 : DFKCNQD1BWP7T port map(CN => FE_PHN393_ml_ms_cntD_n_23, CP => CTS_322, D => FE_PHN500_ml_ms_cntD_n_22, Q => ml_ms_count_debounce(12));
  ml_ms_cntD_count_reg_11 : DFKCNQD1BWP7T port map(CN => FE_PHN393_ml_ms_cntD_n_23, CP => CTS_322, D => ml_ms_cntD_n_21, Q => FE_PHN384_ml_ms_count_debounce_11);
  ml_ms_cntD_g225 : MOAI22D0BWP7T port map(A1 => ml_ms_cntD_n_20, A2 => ml_ms_count_debounce(12), B1 => ml_ms_cntD_n_20, B2 => ml_ms_count_debounce(12), ZN => ml_ms_cntD_n_22);
  ml_ms_cntD_count_reg_10 : DFKCNQD1BWP7T port map(CN => FE_PHN393_ml_ms_cntD_n_23, CP => CTS_322, D => ml_ms_cntD_n_19, Q => FE_PHN379_ml_ms_count_debounce_10);
  ml_ms_cntD_g227 : MOAI22D0BWP7T port map(A1 => ml_ms_cntD_n_18, A2 => ml_ms_count_debounce(11), B1 => ml_ms_cntD_n_18, B2 => ml_ms_count_debounce(11), ZN => ml_ms_cntD_n_21);
  ml_ms_cntD_g228 : IND2D1BWP7T port map(A1 => ml_ms_cntD_n_18, B1 => ml_ms_count_debounce(11), ZN => ml_ms_cntD_n_20);
  ml_ms_cntD_count_reg_9 : DFKCNQD1BWP7T port map(CN => FE_PHN393_ml_ms_cntD_n_23, CP => CTS_322, D => ml_ms_cntD_n_17, Q => ml_ms_count_debounce(9));
  ml_ms_cntD_g230 : MOAI22D0BWP7T port map(A1 => ml_ms_cntD_n_16, A2 => ml_ms_count_debounce(10), B1 => ml_ms_cntD_n_16, B2 => ml_ms_count_debounce(10), ZN => ml_ms_cntD_n_19);
  ml_ms_cntD_g231 : IND2D1BWP7T port map(A1 => ml_ms_cntD_n_16, B1 => ml_ms_count_debounce(10), ZN => ml_ms_cntD_n_18);
  ml_ms_cntD_count_reg_8 : DFKCNQD1BWP7T port map(CN => FE_PHN393_ml_ms_cntD_n_23, CP => CTS_322, D => ml_ms_cntD_n_15, Q => ml_ms_count_debounce(8));
  ml_ms_cntD_g233 : MOAI22D0BWP7T port map(A1 => ml_ms_cntD_n_14, A2 => FE_PHN361_ml_ms_count_debounce_9, B1 => ml_ms_cntD_n_14, B2 => FE_PHN361_ml_ms_count_debounce_9, ZN => ml_ms_cntD_n_17);
  ml_ms_cntD_g234 : IND2D1BWP7T port map(A1 => ml_ms_cntD_n_14, B1 => FE_PHN361_ml_ms_count_debounce_9, ZN => ml_ms_cntD_n_16);
  ml_ms_cntD_count_reg_7 : DFKCNQD1BWP7T port map(CN => FE_PHN393_ml_ms_cntD_n_23, CP => CTS_322, D => FE_PHN498_ml_ms_cntD_n_13, Q => ml_ms_count_debounce(7));
  ml_ms_cntD_g236 : MOAI22D0BWP7T port map(A1 => ml_ms_cntD_n_12, A2 => FE_PHN360_ml_ms_count_debounce_8, B1 => ml_ms_cntD_n_12, B2 => FE_PHN360_ml_ms_count_debounce_8, ZN => ml_ms_cntD_n_15);
  ml_ms_cntD_g237 : IND2D1BWP7T port map(A1 => ml_ms_cntD_n_12, B1 => FE_PHN360_ml_ms_count_debounce_8, ZN => ml_ms_cntD_n_14);
  ml_ms_cntD_count_reg_6 : DFKCNQD1BWP7T port map(CN => FE_PHN393_ml_ms_cntD_n_23, CP => CTS_322, D => ml_ms_cntD_n_11, Q => ml_ms_count_debounce(6));
  ml_ms_cntD_g239 : MOAI22D0BWP7T port map(A1 => FE_PHN489_ml_ms_cntD_n_10, A2 => ml_ms_count_debounce(7), B1 => FE_PHN489_ml_ms_cntD_n_10, B2 => ml_ms_count_debounce(7), ZN => ml_ms_cntD_n_13);
  ml_ms_cntD_g240 : IND2D1BWP7T port map(A1 => FE_PHN489_ml_ms_cntD_n_10, B1 => ml_ms_count_debounce(7), ZN => FE_PHN499_ml_ms_cntD_n_12);
  ml_ms_cntD_count_reg_5 : DFKCNQD1BWP7T port map(CN => FE_PHN393_ml_ms_cntD_n_23, CP => CTS_322, D => FE_PHN491_ml_ms_cntD_n_9, Q => ml_ms_count_debounce(5));
  ml_ms_cntD_g242 : MOAI22D0BWP7T port map(A1 => ml_ms_cntD_n_8, A2 => ml_ms_count_debounce(6), B1 => ml_ms_cntD_n_8, B2 => ml_ms_count_debounce(6), ZN => FE_PHN490_ml_ms_cntD_n_11);
  ml_ms_cntD_g243 : IND2D1BWP7T port map(A1 => ml_ms_cntD_n_8, B1 => ml_ms_count_debounce(6), ZN => ml_ms_cntD_n_10);
  ml_ms_cntD_count_reg_4 : DFKCNQD1BWP7T port map(CN => FE_PHN393_ml_ms_cntD_n_23, CP => CTS_322, D => ml_ms_cntD_n_7, Q => ml_ms_count_debounce(4));
  ml_ms_cntD_g245 : MOAI22D0BWP7T port map(A1 => ml_ms_cntD_n_6, A2 => ml_ms_count_debounce(5), B1 => ml_ms_cntD_n_6, B2 => ml_ms_count_debounce(5), ZN => ml_ms_cntD_n_9);
  ml_ms_cntD_g246 : IND2D1BWP7T port map(A1 => ml_ms_cntD_n_6, B1 => ml_ms_count_debounce(5), ZN => ml_ms_cntD_n_8);
  ml_ms_cntD_count_reg_3 : DFKCNQD1BWP7T port map(CN => FE_PHN393_ml_ms_cntD_n_23, CP => CTS_322, D => ml_ms_cntD_n_5, Q => ml_ms_count_debounce(3));
  ml_ms_cntD_g248 : MOAI22D0BWP7T port map(A1 => ml_ms_cntD_n_4, A2 => FE_PHN375_ml_ms_count_debounce_4, B1 => ml_ms_cntD_n_4, B2 => FE_PHN375_ml_ms_count_debounce_4, ZN => ml_ms_cntD_n_7);
  ml_ms_cntD_g249 : IND2D1BWP7T port map(A1 => ml_ms_cntD_n_4, B1 => FE_PHN375_ml_ms_count_debounce_4, ZN => ml_ms_cntD_n_6);
  ml_ms_cntD_count_reg_2 : DFKCNQD1BWP7T port map(CN => FE_PHN393_ml_ms_cntD_n_23, CP => CTS_322, D => ml_ms_cntD_n_3, Q => ml_ms_cntD_count(2));
  ml_ms_cntD_g251 : MOAI22D0BWP7T port map(A1 => ml_ms_cntD_n_2, A2 => FE_PHN377_ml_ms_count_debounce_3, B1 => ml_ms_cntD_n_2, B2 => FE_PHN377_ml_ms_count_debounce_3, ZN => ml_ms_cntD_n_5);
  ml_ms_cntD_g252 : IND2D1BWP7T port map(A1 => ml_ms_cntD_n_2, B1 => FE_PHN377_ml_ms_count_debounce_3, ZN => ml_ms_cntD_n_4);
  ml_ms_cntD_count_reg_1 : EDFKCND1BWP7T port map(CN => FE_PHN393_ml_ms_cntD_n_23, CP => CTS_322, D => FE_PHN399_ml_ms_cntD_count_1, E => ml_ms_cntD_count(0), Q => UNCONNECTED17, QN => ml_ms_cntD_count(1));
  ml_ms_cntD_g254 : MOAI22D0BWP7T port map(A1 => ml_ms_cntD_n_1, A2 => FE_PHN356_ml_ms_cntD_count_2, B1 => ml_ms_cntD_n_1, B2 => FE_PHN356_ml_ms_cntD_count_2, ZN => ml_ms_cntD_n_3);
  ml_ms_cntD_g255 : IND2D1BWP7T port map(A1 => ml_ms_cntD_n_1, B1 => FE_PHN356_ml_ms_cntD_count_2, ZN => ml_ms_cntD_n_2);
  ml_ms_cntD_g257 : IND2D1BWP7T port map(A1 => FE_PHN399_ml_ms_cntD_count_1, B1 => ml_ms_cntD_count(0), ZN => ml_ms_cntD_n_1);
  ml_ms_cntD_count_reg_0 : DFKCND1BWP7T port map(CN => FE_PHN397_ml_ms_cntD_n_0, CP => CTS_322, D => FE_PHN393_ml_ms_cntD_n_23, Q => FE_PHN357_ml_ms_cntD_count_0, QN => ml_ms_cntD_n_0);
  tie_1_cell : TIEHBWP7T port map(Z => logic_1_1_net);

end routed;
