configuration e_counter_behav_cfg of e_counter is
   for behav
   end for;
end e_counter_behav_cfg;
