configuration y_behaviour_y_cfg of y is
   for behaviour_y
   end for;
end y_behaviour_y_cfg;
