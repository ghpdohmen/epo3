library IEEE;
use IEEE.std_logic_1164.ALL;

entity vgatest_tb is
end vgatest_tb;

