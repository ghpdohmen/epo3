configuration mouse_tb_behav_cfg2 of mouse_tb is
   for behav
      for all: mouse use configuration work.mouse_synthesised_cfg;
      end for;
   end for;
end mouse_tb_behav_cfg2;
