configuration vgadriver_behaviour_cfg of vgadriver is
   for behaviour
   end for;
end vgadriver_behaviour_cfg;
