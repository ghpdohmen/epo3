configuration graphic_toplvl_tb_behaviour_cfg of graphic_toplvl_tb is
   for behaviour
      for all: graphic_toplvl use configuration work.graphic_toplvl_behaviour_cfg;
      end for;
   end for;
end graphic_toplvl_tb_behaviour_cfg;
