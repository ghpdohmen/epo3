configuration mouse_synthesised_cfg of mouse is
   for synthesised
      -- skipping invd1bwp7t because it is not a local entity
      -- skipping buffd4bwp7t because it is not a local entity
      -- skipping nr2xd0bwp7t because it is not a local entity
      -- skipping dfqd1bwp7t because it is not a local entity
      -- skipping dfd1bwp7t because it is not a local entity
      -- skipping inr2d0bwp7t because it is not a local entity
      -- skipping ind3d1bwp7t because it is not a local entity
      -- skipping oai221d0bwp7t because it is not a local entity
      -- skipping an2d0bwp7t because it is not a local entity
      -- skipping an2d1bwp7t because it is not a local entity
      -- skipping ind2d1bwp7t because it is not a local entity
      -- skipping an2d4bwp7t because it is not a local entity
      -- skipping maoi22d0bwp7t because it is not a local entity
      -- skipping an3d1bwp7t because it is not a local entity
      -- skipping nd2d1bwp7t because it is not a local entity
      -- skipping nd2d0bwp7t because it is not a local entity
      -- skipping inr3d0bwp7t because it is not a local entity
      -- skipping moai22d0bwp7t because it is not a local entity
      -- skipping dfqd0bwp7t because it is not a local entity
      -- skipping oai21d0bwp7t because it is not a local entity
      -- skipping aoi21d0bwp7t because it is not a local entity
      -- skipping aoi222d0bwp7t because it is not a local entity
      -- skipping oai211d1bwp7t because it is not a local entity
      -- skipping oai31d0bwp7t because it is not a local entity
      -- skipping aoi32d1bwp7t because it is not a local entity
      -- skipping ao21d0bwp7t because it is not a local entity
      -- skipping ioa21d1bwp7t because it is not a local entity
      -- skipping iao21d0bwp7t because it is not a local entity
      -- skipping aoi33d1bwp7t because it is not a local entity
      -- skipping nr2d1bwp7t because it is not a local entity
      -- skipping invd0bwp7t because it is not a local entity
      -- skipping or2d1bwp7t because it is not a local entity
      -- skipping inr2d1bwp7t because it is not a local entity
      -- skipping edfqd0bwp7t because it is not a local entity
      -- skipping aoi22d0bwp7t because it is not a local entity
      -- skipping dfkcnqd1bwp7t because it is not a local entity
      -- skipping ckxor2d0bwp7t because it is not a local entity
      -- skipping edfkcnqd1bwp7t because it is not a local entity
      -- skipping lhqd1bwp7t because it is not a local entity
      -- skipping ioa21d0bwp7t because it is not a local entity
      -- skipping aoi221d0bwp7t because it is not a local entity
      -- skipping nd4d0bwp7t because it is not a local entity
      -- skipping cknd1bwp7t because it is not a local entity
      -- skipping nd3d0bwp7t because it is not a local entity
      -- skipping nr2d0bwp7t because it is not a local entity
      -- skipping inr2xd0bwp7t because it is not a local entity
      -- skipping cknd2d1bwp7t because it is not a local entity
      -- skipping dfkcnd1bwp7t because it is not a local entity
      -- skipping ao221d0bwp7t because it is not a local entity
      -- skipping ao22d0bwp7t because it is not a local entity
      -- skipping nd2d4bwp7t because it is not a local entity
   end for;
end mouse_synthesised_cfg;
