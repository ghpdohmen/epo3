configuration flipflop_behav_cfg of flipflop is
   for behav
   end for;
end flipflop_behav_cfg;
