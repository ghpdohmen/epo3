configuration counter25mhz_synthesised_cfg of counter25mhz is
   for synthesised
      -- skipping ind2d1bwp7t because it is not a local entity
      -- skipping dfkcnqd1bwp7t because it is not a local entity
      -- skipping moai22d0bwp7t because it is not a local entity
      -- skipping nd2d1bwp7t because it is not a local entity
      -- skipping buffd4bwp7t because it is not a local entity
      -- skipping invd1bwp7t because it is not a local entity
      -- skipping xnr2d1bwp7t because it is not a local entity
      -- skipping invd4bwp7t because it is not a local entity
      -- skipping dfkcnd1bwp7t because it is not a local entity
      -- skipping dfkcnd0bwp7t because it is not a local entity
   end for;
end counter25mhz_synthesised_cfg;
