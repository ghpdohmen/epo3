configuration shiftregister_9bit_tb_behav_cfg of shiftregister_9bit_tb is
   for behav
      for all: shiftregister_9bit use configuration work.shiftregister_9bit_behav_cfg;
      end for;
   end for;
end shiftregister_9bit_tb_behav_cfg;
