configuration shiftregister_11bit_tb_behaviour_cfg of shiftregister_11bit_tb is
   for behaviour
      for all: shiftregister_11bit use configuration work.shiftregister_11bit_behav_cfg;
      end for;
   end for;
end shiftregister_11bit_tb_behaviour_cfg;
