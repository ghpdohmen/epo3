configuration counter25mhz_behav_cfg of counter25mhz is
   for behav
   end for;
end counter25mhz_behav_cfg;
