configuration x_behaviour_x_cfg of x is
   for behaviour_x
   end for;
end x_behaviour_x_cfg;
