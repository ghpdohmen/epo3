configuration submod_vcount_behaviour_cfg of submod_vcount is
   for behaviour
   end for;
end submod_vcount_behaviour_cfg;
