configuration shiftregister_9bit_synthesised_cfg of shiftregister_9bit is
   for synthesised
      -- skipping dfqd1bwp7t because it is not a local entity
      -- skipping ao222d0bwp7t because it is not a local entity
      -- skipping ao22d0bwp7t because it is not a local entity
      -- skipping nr2d1bwp7t because it is not a local entity
      -- skipping an2d1bwp7t because it is not a local entity
      -- skipping cknd1bwp7t because it is not a local entity
      -- skipping invd4bwp7t because it is not a local entity
      -- skipping dfd0bwp7t because it is not a local entity
   end for;
end shiftregister_9bit_synthesised_cfg;
