configuration pixel_behav_cfg of pixel is
   for behav
