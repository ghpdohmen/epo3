configuration submod_ecount_behaviour_cfg of submod_ecount is
   for behaviour
   end for;
end submod_ecount_behaviour_cfg;
