configuration sendfsm_behav_cfg of sendfsm is
   for behav
   end for;
end sendfsm_behav_cfg;
