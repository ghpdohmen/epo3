configuration timebase_synthesised_cfg of timebase is
   for synthesised
      -- skipping ao32d1bwp7t because it is not a local entity
      -- skipping oai21d0bwp7t because it is not a local entity
      -- skipping moai22d0bwp7t because it is not a local entity
      -- skipping invd0bwp7t because it is not a local entity
      -- skipping oai22d0bwp7t because it is not a local entity
      -- skipping nr2xd0bwp7t because it is not a local entity
      -- skipping iao21d0bwp7t because it is not a local entity
      -- skipping cknd2d0bwp7t because it is not a local entity
      -- skipping ind3d1bwp7t because it is not a local entity
      -- skipping mux2d0bwp7t because it is not a local entity
      -- skipping inr2d0bwp7t because it is not a local entity
      -- skipping invd4bwp7t because it is not a local entity
      -- skipping dfd0bwp7t because it is not a local entity
   end for;
end timebase_synthesised_cfg;
