configuration shiftregister_11bit_tb_behav_cfg2 of shiftregister_11bit_tb is
   for behav
      for all: shiftregister_11bit use configuration work.shiftregister_11bit_synthesised_cfg;
      end for;
   end for;
end shiftregister_11bit_tb_behav_cfg2;
