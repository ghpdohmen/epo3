library IEEE;
use IEEE.std_logic_1164.ALL;

entity buffer is
   port(input  : in  std_logic;
        clk    : in  std_logic;
        output : out std_logic);
end buffer;

