configuration color_behaviour_color_cfg of color is
   for behaviour_color
   end for;
end color_behaviour_color_cfg;
