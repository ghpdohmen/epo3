configuration mouse_tb_behav_cfg_routed of mouse_tb is
   for behav
      for all: mouse use configuration work.mouse_routed_cfg;
      end for;
   end for;
end mouse_tb_behav_cfg_routed;
