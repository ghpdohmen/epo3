
library ieee;
use ieee.std_logic_1164.all;
--library tcb018gbwp7t;
--use tcb018gbwp7t.all;

architecture synthesised of pixel is

  component mouse_timer
    port(clk       : in  std_logic;
         reset     : in  std_logic;
         count_out : out std_logic_vector(21 downto 0));
  end component;

  component BUFFD4BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component LHQD1BWP7T
    port(E, D : in std_logic; Q : out std_logic);
  end component;

  component MOAI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component ND4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component AN4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component AOI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AN2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component INR2D1BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component NR2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component AN2D4BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component NR2XD0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component NR2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component ND2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component CKND2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component INVD0BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component IND2D1BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component INVD2BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component XNR2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component INR2D0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component ND2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component CKND1BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component FA1D0BWP7T
    port(A, B, CI : in std_logic; CO, S : out std_logic);
  end component;

  component IND2D0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component INVD1BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component HA1D0BWP7T
    port(A, B : in std_logic; CO, S : out std_logic);
  end component;

  component DFQD1BWP7T
    port(CP, D : in std_logic; Q : out std_logic);
  end component;

  component DFQD0BWP7T
    port(CP, D : in std_logic; Q : out std_logic);
  end component;

  component AO221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; Z : out std_logic);
  end component;

  component AO22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component INR2XD0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component OAI211D1BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component AOI211XD0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component AO32D1BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component OAI21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component AOI21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component CKAN2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component AN4D1BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component NR4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component OA21D0BWP7T
    port(A1, A2, B : in std_logic; Z : out std_logic);
  end component;

  component MAOI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component DFD1BWP7T
    port(CP, D : in std_logic; Q, QN : out std_logic);
  end component;

  component DFD0BWP7T
    port(CP, D : in std_logic; Q, QN : out std_logic);
  end component;

  component OR2D4BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component OAI221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; ZN : out std_logic);
  end component;

  component IND3D1BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component IAO21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component IOA21D1BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component OA31D1BWP7T
    port(A1, A2, A3, B : in std_logic; Z : out std_logic);
  end component;

  component OA22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component AO211D0BWP7T
    port(A1, A2, B, C : in std_logic; Z : out std_logic);
  end component;

  component AN2D0BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component OR2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component NR3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component AO21D0BWP7T
    port(A1, A2, B : in std_logic; Z : out std_logic);
  end component;

  component OAI31D0BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component AN3D0BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component OR4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component OA31D0BWP7T
    port(A1, A2, A3, B : in std_logic; Z : out std_logic);
  end component;

  component ND3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component AOI32D1BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OA211D0BWP7T
    port(A1, A2, B, C : in std_logic; Z : out std_logic);
  end component;

  component AO33D0BWP7T
    port(A1, A2, A3, B1, B2, B3 : in std_logic; Z : out std_logic);
  end component;

  component OAI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AOI222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; ZN : out std_logic);
  end component;

  component OR4D1BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component DFKCND1BWP7T
    port(CP, CN, D : in std_logic; Q, QN : out std_logic);
  end component;

  component DFXD1BWP7T
    port(CP, DA, DB, SA : in std_logic; Q, QN : out std_logic);
  end component;

  component EDFQD1BWP7T
    port(CP, D, E : in std_logic; Q : out std_logic);
  end component;

  component EDFQD0BWP7T
    port(CP, D, E : in std_logic; Q : out std_logic);
  end component;

  component EDFKCNQD1BWP7T
    port(CP, CN, D, E : in std_logic; Q : out std_logic);
  end component;

  component DFKCNQD1BWP7T
    port(CP, CN, D : in std_logic; Q : out std_logic);
  end component;

  component CKXOR2D0BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component CKXOR2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component DFKSND1BWP7T
    port(CP, D, SN : in std_logic; Q, QN : out std_logic);
  end component;

  component OR3D1BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component INR3D0BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component DFXQD1BWP7T
    port(CP, DA, DB, SA : in std_logic; Q : out std_logic);
  end component;

  component ND2D4BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component EDFKCND1BWP7T
    port(CP, CN, D, E : in std_logic; Q, QN : out std_logic);
  end component;

  component INR4D0BWP7T
    port(A1, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component OAI32D1BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component IND4D0BWP7T
    port(A1, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component AOI31D0BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component OR3D4BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component IINR4D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component MUX2ND0BWP7T
    port(I0, I1, S : in std_logic; ZN : out std_logic);
  end component;

  component MUX2D1BWP7T
    port(I0, I1, S : in std_logic; Z : out std_logic);
  end component;

  component LNQD1BWP7T
    port(EN, D : in std_logic; Q : out std_logic);
  end component;

  component AOI211D1BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component OAI222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; ZN : out std_logic);
  end component;

  component AOI221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; ZN : out std_logic);
  end component;

  component OAI33D1BWP7T
    port(A1, A2, A3, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component AOI33D1BWP7T
    port(A1, A2, A3, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component DFKCNQD2BWP7T
    port(CP, CN, D : in std_logic; Q : out std_logic);
  end component;

  component OAI32D0BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  signal gl_sig_rom : std_logic_vector(1 downto 0);
  signal gl_sig_e : std_logic_vector(9 downto 0);
  signal gl_rom_rom_776 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_779 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_385 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_389 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_977 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_981 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_980 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_982 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_384 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_387 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_978 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_979 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_976 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_983 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_712 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_713 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_956 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_958 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_882 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_887 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_706 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_711 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_985 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_989 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_988 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_990 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_378 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_383 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_986 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_987 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_984 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_991 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_708 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_710 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_380 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_382 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_994 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_999 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_993 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_997 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_880 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_883 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_381 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_379 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_996 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_998 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_376 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_377 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_992 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_995 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1022 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1023 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_709 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_707 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1020 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1018 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_362 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_367 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_704 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_705 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1017 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1021 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1016 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1019 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_361 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_365 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1006 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1007 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1004 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1002 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_364 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_366 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_360 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_363 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1001 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1005 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1000 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1003 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_974 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_975 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_957 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_955 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_972 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_970 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_370 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_375 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_969 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_973 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_854 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_855 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_968 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_971 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_372 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_374 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_794 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_799 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_966 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_967 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_373 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_371 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_964 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_962 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_852 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_850 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_961 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_965 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_960 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_963 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_368 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_369 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_953 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_793 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_797 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_796 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_798 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_338 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_343 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_954 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_340 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_342 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_952 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_959 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_792 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_795 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_937 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_941 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_341 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_339 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_940 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_942 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_938 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_939 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_336 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_337 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_936 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_943 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_926 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_927 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_849 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_853 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_924 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_922 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_346 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_351 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_921 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_925 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_801 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_805 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_920 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_923 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_348 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_350 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_848 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_851 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_930 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_935 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_929 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_933 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_349 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_347 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_932 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_934 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_344 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_345 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_928 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_931 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_804 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_806 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_945 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_949 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_948 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_950 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_354 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_359 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_802 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_807 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_946 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_947 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_356 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_358 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_944 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_951 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_914 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_919 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_800 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_803 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_357 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_355 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_913 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_917 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_352 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_353 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_916 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_915 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_912 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_918 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_905 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_909 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_908 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_910 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_329 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_333 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_906 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_911 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_904 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_907 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_332 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_334 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_817 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_821 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_898 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_903 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_890 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_895 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_330 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_331 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_897 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_901 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_820 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_822 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_328 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_335 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_900 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_902 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_896 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_899 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_892 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_894 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_702 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_703 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_322 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_327 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_700 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_698 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_818 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_819 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_697 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_701 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_696 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_699 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_324 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_326 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_325 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_323 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_686 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_687 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_816 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_823 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_684 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_682 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_320 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_321 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_681 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_685 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_680 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_683 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_893 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_891 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_690 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_695 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_692 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_694 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_126 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_127 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_693 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_691 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_688 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_689 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_124 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_122 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_662 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_663 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_786 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_791 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_660 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_658 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_785 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_789 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_121 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_125 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_120 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_123 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_657 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_661 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_656 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_659 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_666 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_671 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_888 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_889 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_788 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_787 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_665 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_669 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_106 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_111 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_105 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_109 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_668 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_667 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_664 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_670 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_678 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_679 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_784 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_790 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_108 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_107 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_676 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_674 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_104 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_110 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_673 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_677 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_672 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_675 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_654 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_655 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_652 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_650 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_874 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_879 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_114 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_119 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_649 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_653 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_116 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_118 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_648 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_651 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_825 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_829 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_828 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_830 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_642 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_647 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_117 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_115 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_641 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_645 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_644 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_646 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_640 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_643 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_569 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_573 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_112 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_113 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_873 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_877 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_82 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_87 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_572 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_574 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_826 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_827 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_570 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_571 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_84 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_86 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_568 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_575 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_824 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_831 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_85 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_83 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_554 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_559 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_553 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_557 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_556 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_558 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_80 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_81 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_552 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_555 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_876 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_875 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_566 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_567 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_564 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_562 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_90 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_95 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_810 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_815 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_561 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_565 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_92 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_94 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_560 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_563 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_534 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_535 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_93 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_91 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_532 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_530 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_809 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_813 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_529 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_533 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_528 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_531 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_88 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_89 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_542 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_543 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_872 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_878 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_812 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_811 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_102 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_103 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_540 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_538 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_100 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_98 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_537 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_541 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_536 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_539 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_550 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_551 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_808 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_814 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_97 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_101 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_548 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_546 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_96 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_99 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_545 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_549 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_544 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_547 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_526 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_527 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_524 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_522 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_74 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_79 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_842 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_847 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_521 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_525 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_778 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_783 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_520 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_523 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_73 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_77 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_513 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_517 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_76 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_75 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_516 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_518 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_72 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_78 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_514 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_519 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_512 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_515 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_777 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_781 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_66 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_71 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_780 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_782 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_498 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_503 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_497 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_501 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_841 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_845 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_68 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_70 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_500 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_502 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_496 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_499 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_69 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_67 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1008 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1011 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_465 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_469 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_468 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_470 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_64 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_65 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_466 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_471 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_464 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_467 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_844 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_843 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_474 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_479 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_770 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_775 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_476 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_478 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_217 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_221 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_477 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_475 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_472 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_473 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_220 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_222 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_769 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_773 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_486 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_487 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_484 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_482 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_218 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_219 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_481 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_485 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_480 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_483 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_216 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_223 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_506 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_511 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_840 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_846 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_772 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_774 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_225 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_229 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_508 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_510 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_768 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_771 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_509 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_507 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_228 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_230 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_504 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_505 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_489 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_493 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_226 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_227 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_492 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_494 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1012 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1014 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_490 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_495 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_224 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_231 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_488 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_491 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_834 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_839 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_458 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_463 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_457 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_461 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_242 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_247 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_460 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_462 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_456 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_459 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_241 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_245 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_449 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_453 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_244 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_246 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_452 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_454 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_450 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_455 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_240 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_243 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_448 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_451 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_833 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_837 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_442 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_447 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_214 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_215 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_444 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_446 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_212 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_210 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_445 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_443 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_440 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_441 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_426 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_431 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_209 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_213 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_425 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_429 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_428 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_430 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_424 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_427 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_208 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_211 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_836 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_835 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_410 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_415 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_409 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_413 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_254 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_255 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_412 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_414 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_252 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_250 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_408 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_411 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_832 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_838 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_422 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_423 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_249 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_253 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_420 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_418 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_417 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_421 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_416 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_419 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_248 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_251 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_433 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_437 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_436 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_438 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_233 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_237 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_434 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_439 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_236 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_238 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_432 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_435 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_402 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_407 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_234 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_235 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_401 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_405 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_404 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_406 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_232 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_239 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_400 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_403 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_393 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_397 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_396 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_398 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_201 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_205 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_394 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_399 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_204 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_206 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_392 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_395 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_390 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_391 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_634 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_639 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_388 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_386 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_202 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_203 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_200 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_207 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_193 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_197 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_196 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_198 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_636 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_638 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_194 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_195 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_192 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_199 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_637 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_635 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_318 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_319 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_316 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_314 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_313 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_317 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_312 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_315 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_302 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_303 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_632 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_633 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_300 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_298 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_297 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_301 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_296 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_299 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_281 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_285 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_284 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_286 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_282 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_283 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_617 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_621 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_280 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_287 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_620 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_622 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_289 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_293 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_292 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_294 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_290 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_291 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_288 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_295 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_618 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_619 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_310 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_311 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_308 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_306 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_305 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_309 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_304 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_307 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_274 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_279 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_273 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_277 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_276 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_278 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_272 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_275 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_616 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_623 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_270 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_271 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_266 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_268 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_265 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_269 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_264 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_267 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_602 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_607 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_258 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_263 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_257 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_261 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_260 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_262 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_256 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_259 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_604 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_606 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_605 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_603 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_190 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_191 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_188 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_186 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_185 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_189 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_184 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_187 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_600 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_601 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_169 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_173 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_172 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_174 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_170 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_171 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_168 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_175 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_154 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_159 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_610 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_615 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_156 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_158 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_157 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_155 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_152 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_153 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_609 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_613 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_166 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_167 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_164 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_162 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_161 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_165 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_160 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_163 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_612 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_611 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_178 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_183 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_608 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_614 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_180 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_182 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_181 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_179 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_176 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_177 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_146 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_151 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_148 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_150 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_149 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_147 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_144 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_145 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_138 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_143 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_625 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_629 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_140 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_142 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_141 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_139 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_136 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_137 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_130 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_135 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_628 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_630 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_129 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_133 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_132 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_134 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_128 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_131 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_626 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_627 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_58 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_63 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_57 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_61 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_60 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_62 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_56 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_59 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_624 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_631 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_46 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_47 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_44 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_42 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_41 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_45 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_40 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_43 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1013 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_594 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_599 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_50 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_55 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_52 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_54 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_53 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_51 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_48 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_49 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_593 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_597 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_17 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_21 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_20 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_22 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_18 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_19 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_16 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_23 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_596 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_598 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_26 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_31 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_25 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_29 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_28 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_27 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_592 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_595 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_24 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_30 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_34 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_39 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_36 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_38 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_37 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_35 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_33 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_32 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_9 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_13 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_14 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_15 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_12 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_10 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_11 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_586 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_591 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_8 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_2 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_7 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_5 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_588 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_590 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_4 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_6 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_0 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_3 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_589 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_587 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_584 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_585 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_578 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_583 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_580 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_582 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_862 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_863 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_860 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_858 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_857 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_861 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_856 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_859 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_870 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_871 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_868 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_866 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_581 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_579 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_865 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_869 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_864 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_867 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_886 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_884 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_576 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_577 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_881 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_885 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_754 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_759 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_753 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_757 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_756 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_755 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_752 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_758 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_722 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_727 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_724 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_726 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1009 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_725 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_723 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_720 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_721 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_730 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_735 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_729 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_733 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_761 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_765 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_732 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_731 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_764 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_766 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_762 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_767 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_760 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_763 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_728 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_734 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_746 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_751 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_748 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_750 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_749 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_747 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_744 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_745 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_738 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_743 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_740 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_742 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_741 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_739 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_736 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_737 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_714 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_719 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_716 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_718 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_717 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_715 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1010 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1015 : std_logic_vector(1 downto 0);
  signal gl_sig_ram : std_logic_vector(2 downto 0);
  signal gl_ram_ram_96 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_97 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_98 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_99 : std_logic_vector(2 downto 0);
  signal gl_sig_y : std_logic_vector(3 downto 0);
  signal gl_ram_ram_80 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_83 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_41 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_42 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_78 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_79 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_62 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_63 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_60 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_61 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_44 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_45 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_57 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_58 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_40 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_43 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_56 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_59 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_72 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_75 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_54 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_55 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_49 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_50 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_52 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_53 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_38 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_39 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_48 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_51 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_33 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_34 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_30 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_31 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_24 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_27 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_36 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_37 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_28 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_29 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_94 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_95 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_25 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_26 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_32 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_35 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_14 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_15 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_12 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_13 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_66 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_67 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_10 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_11 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_88 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_91 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_8 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_9 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_46 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_47 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_92 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_93 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_89 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_90 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_22 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_23 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_16 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_19 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_20 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_21 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_17 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_18 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_70 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_71 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_6 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_7 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_1 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_2 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_4 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_5 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_0 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_3 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_86 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_87 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_65 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_68 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_69 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_84 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_85 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_81 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_82 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_64 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_73 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_74 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_76 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_77 : std_logic_vector(2 downto 0);
  signal gl_sig_x : std_logic_vector(3 downto 0);
  signal gl_ram_ram_position : std_logic_vector(6 downto 0);
  signal gl_ram_x_grid : std_logic_vector(6 downto 0);
  signal gl_ram_y_grid : std_logic_vector(6 downto 0);
  signal sig_output_color : std_logic_vector(2 downto 0);
  signal sig_logic_y : std_logic_vector(3 downto 0);
  signal sig_logic_x : std_logic_vector(3 downto 0);
  signal ml_mouseX : std_logic_vector(2 downto 0);
  signal ml_buttons_mouse : std_logic_vector(4 downto 0);
  signal ml_ms_timer_count : std_logic_vector(21 downto 0);
  signal ml_ms_sfsm_state : std_logic_vector(3 downto 0);
  signal ml_ms_sr_new_new_data : std_logic_vector(8 downto 0);
  signal ml_ms_count25M : std_logic_vector(12 downto 0);
  signal ml_ms_data_sr_11bit : std_logic_vector(10 downto 0);
  signal ml_ms_mouse_x : std_logic_vector(2 downto 0);
  signal ml_ms_mouse_y : std_logic_vector(2 downto 0);
  signal ml_ms_mfsm_state : std_logic_vector(4 downto 0);
  signal ml_ms_btns : std_logic_vector(4 downto 0);
  signal ml_ms_count15k : std_logic_vector(3 downto 0);
  signal ml_il_y1_locy : std_logic_vector(3 downto 0);
  signal ml_il_y1_input_register : std_logic_vector(3 downto 0);
  signal ml_ms_cnt_count : std_logic_vector(12 downto 0);
  signal ml_il_color1_state : std_logic_vector(2 downto 0);
  signal ml_il_color1_state_hs : std_logic_vector(1 downto 0);
  signal ml_il_x1_input_register : std_logic_vector(3 downto 0);
  signal gl_vgd_horizontal : std_logic_vector(9 downto 0);
  signal gl_vgd_vertical : std_logic_vector(9 downto 0);
  signal gl_vgd_horizontal_counter : std_logic_vector(9 downto 0);
  signal gl_vgd_vertical_counter : std_logic_vector(9 downto 0);
  signal gl_gr_lg_local_y : std_logic_vector(3 downto 0);
  signal gl_gr_lg_local_x : std_logic_vector(3 downto 0);
  signal gl_gr_lg_countdown_case : std_logic_vector(10 downto 0);
  signal gl_gr_lg_le_new_count_e : std_logic_vector(9 downto 0);
  signal gl_gr_lg_le_x_old : std_logic_vector(3 downto 0);
  signal gl_gr_lg_le_y_old : std_logic_vector(3 downto 0);
  signal ml_ms_ed_state : std_logic_vector(1 downto 0);
  signal ml_ms_count_debounce : std_logic_vector(12 downto 0);
  signal ml_ms_cntD_count : std_logic_vector(12 downto 0);
  signal UNCONNECTED, UNCONNECTED0, UNCONNECTED1, UNCONNECTED2, gl_gr_lg_lcountdown_l_edge_reg1 : std_logic;
  signal gl_gr_lg_lcountdown_l_edge_reg2, gl_gr_lg_lcountdown_n_0, gl_gr_lg_lcountdown_n_1, gl_gr_lg_lcountdown_n_2, gl_gr_lg_lcountdown_n_3 : std_logic;
  signal gl_gr_lg_lcountdown_n_4, gl_gr_lg_lcountdown_n_5, gl_gr_lg_lcountdown_n_6, gl_gr_lg_lcountdown_n_7, gl_gr_lg_lcountdown_n_8 : std_logic;
  signal gl_gr_lg_lcountdown_n_9, gl_gr_lg_lcountdown_n_10, gl_gr_lg_lcountdown_n_11, gl_gr_lg_lcountdown_n_12, gl_gr_lg_lcountdown_n_13 : std_logic;
  signal gl_gr_lg_lcountdown_n_14, gl_gr_lg_lcountdown_n_15, gl_gr_lg_lcountdown_n_16, gl_gr_lg_lcountdown_n_17, gl_gr_lg_lcountdown_n_18 : std_logic;
  signal gl_gr_lg_lcountdown_n_19, gl_gr_lg_lcountdown_n_20, gl_gr_lg_lcountdown_n_21, gl_gr_lg_lcountdown_n_22, gl_gr_lg_lcountdown_n_23 : std_logic;
  signal gl_gr_lg_lcountdown_n_24, gl_gr_lg_lcountdown_n_25, gl_gr_lg_lcountdown_n_26, gl_gr_lg_lcountdown_n_27, gl_gr_lg_lcountdown_n_28 : std_logic;
  signal gl_gr_lg_lcountdown_n_29, gl_gr_lg_lcountdown_n_30, gl_gr_lg_lcountdown_n_31, gl_gr_lg_lcountdown_n_32, gl_gr_lg_lcountdown_n_33 : std_logic;
  signal gl_gr_lg_lcountdown_n_34, gl_gr_lg_lcountdown_n_35, gl_gr_lg_lcountdown_n_36, gl_gr_lg_lcountdown_n_37, gl_gr_lg_lcountdown_n_38 : std_logic;
  signal gl_gr_lg_lcountdown_sig_edge_fall, gl_gr_lg_le_n_0, gl_gr_lg_le_n_1, gl_gr_lg_le_n_2, gl_gr_lg_le_n_3 : std_logic;
  signal gl_gr_lg_le_n_4, gl_gr_lg_le_n_5, gl_gr_lg_le_n_6, gl_gr_lg_le_n_7, gl_gr_lg_le_n_8 : std_logic;
  signal gl_gr_lg_le_n_9, gl_gr_lg_le_n_10, gl_gr_lg_le_n_11, gl_gr_lg_le_n_12, gl_gr_lg_le_n_13 : std_logic;
  signal gl_gr_lg_le_n_14, gl_gr_lg_le_n_15, gl_gr_lg_le_n_16, gl_gr_lg_le_n_17, gl_gr_lg_le_n_18 : std_logic;
  signal gl_gr_lg_le_n_19, gl_gr_lg_le_n_20, gl_gr_lg_le_n_21, gl_gr_lg_le_n_22, gl_gr_lg_le_n_23 : std_logic;
  signal gl_gr_lg_le_n_24, gl_gr_lg_le_n_25, gl_gr_lg_le_n_26, gl_gr_lg_le_n_27, gl_gr_lg_le_n_28 : std_logic;
  signal gl_gr_lg_le_n_29, gl_gr_lg_le_n_30, gl_gr_lg_le_n_31, gl_gr_lg_le_n_32, gl_gr_lg_le_n_33 : std_logic;
  signal gl_gr_lg_le_n_34, gl_gr_lg_le_n_35, gl_gr_lg_le_n_36, gl_gr_lg_le_n_37, gl_gr_lg_le_n_38 : std_logic;
  signal gl_gr_lg_le_n_39, gl_gr_lg_le_n_40, gl_gr_lg_le_n_41, gl_gr_lg_le_n_42, gl_gr_lg_lh_l_edge_n_0 : std_logic;
  signal gl_gr_lg_lh_l_edge_reg1, gl_gr_lg_lh_l_edge_reg2, gl_gr_lg_lh_n_1, gl_gr_lg_lh_n_2, gl_gr_lg_lh_n_3 : std_logic;
  signal gl_gr_lg_lh_n_4, gl_gr_lg_lh_n_5, gl_gr_lg_lh_n_6, gl_gr_lg_lh_n_8, gl_gr_lg_lh_n_10 : std_logic;
  signal gl_gr_lg_lh_n_11, gl_gr_lg_lh_n_12, gl_gr_lg_lh_n_13, gl_gr_lg_lh_n_14, gl_gr_lg_lh_n_15 : std_logic;
  signal gl_gr_lg_lh_n_19, gl_gr_lg_lh_sig_edges, gl_gr_lg_lv_l_edge_n_0, gl_gr_lg_lv_l_edge_reg1, gl_gr_lg_lv_l_edge_reg2 : std_logic;
  signal gl_gr_lg_lv_n_1, gl_gr_lg_lv_n_2, gl_gr_lg_lv_n_3, gl_gr_lg_lv_n_4, gl_gr_lg_lv_n_5 : std_logic;
  signal gl_gr_lg_lv_n_6, gl_gr_lg_lv_n_8, gl_gr_lg_lv_n_10, gl_gr_lg_lv_n_11, gl_gr_lg_lv_n_12 : std_logic;
  signal gl_gr_lg_lv_n_13, gl_gr_lg_lv_n_14, gl_gr_lg_lv_n_15, gl_gr_lg_lv_n_19, gl_gr_lg_lv_sig_edges : std_logic;
  signal gl_gr_lg_n_0, gl_gr_lg_n_1, gl_gr_lg_n_2, gl_gr_lg_n_3, gl_gr_lg_n_4 : std_logic;
  signal gl_gr_lg_n_6, gl_gr_lg_n_7, gl_gr_lg_n_8, gl_gr_lg_n_9, gl_gr_lg_n_10 : std_logic;
  signal gl_gr_lg_n_11, gl_gr_lg_n_12, gl_gr_lg_n_13, gl_gr_lg_n_14, gl_gr_lg_n_15 : std_logic;
  signal gl_gr_lg_n_16, gl_gr_lg_n_17, gl_gr_lg_n_18, gl_gr_lg_n_19, gl_gr_lg_n_20 : std_logic;
  signal gl_gr_lg_n_21, gl_gr_lg_n_22, gl_gr_lg_n_23, gl_gr_lg_n_24, gl_gr_lg_n_25 : std_logic;
  signal gl_gr_lg_n_26, gl_gr_lg_n_27, gl_gr_lg_n_28, gl_gr_lg_n_29, gl_gr_lg_n_30 : std_logic;
  signal gl_gr_lg_n_31, gl_gr_lg_n_32, gl_gr_lg_n_33, gl_gr_lg_n_34, gl_gr_lg_n_35 : std_logic;
  signal gl_gr_lg_n_36, gl_gr_lg_n_37, gl_gr_lg_n_38, gl_gr_lg_n_39, gl_gr_lg_n_40 : std_logic;
  signal gl_gr_lg_n_41, gl_gr_lg_n_42, gl_gr_lg_n_43, gl_gr_lg_n_44, gl_gr_lg_n_45 : std_logic;
  signal gl_gr_lg_n_47, gl_gr_lg_n_48, gl_gr_lg_n_49, gl_gr_lg_n_50, gl_gr_lg_n_51 : std_logic;
  signal gl_gr_lg_n_52, gl_gr_lg_n_53, gl_gr_lg_n_54, gl_gr_lg_n_55, gl_gr_lg_n_56 : std_logic;
  signal gl_gr_lg_n_57, gl_gr_lg_n_58, gl_gr_lg_n_59, gl_gr_lg_n_60, gl_gr_lg_n_61 : std_logic;
  signal gl_gr_lg_n_62, gl_gr_lg_n_63, gl_gr_lg_n_64, gl_gr_lg_n_65, gl_gr_lg_n_66 : std_logic;
  signal gl_gr_lg_n_67, gl_gr_lg_n_68, gl_gr_lg_n_69, gl_gr_lg_n_70, gl_gr_lg_n_71 : std_logic;
  signal gl_gr_lg_n_72, gl_gr_lg_n_73, gl_gr_lg_n_74, gl_gr_lg_n_75, gl_gr_lg_n_76 : std_logic;
  signal gl_gr_lg_n_77, gl_gr_lg_n_78, gl_gr_lg_n_79, gl_gr_lg_n_80, gl_gr_lg_n_81 : std_logic;
  signal gl_gr_lg_n_82, gl_gr_lg_n_83, gl_gr_lg_n_85, gl_gr_lg_n_86, gl_gr_lg_n_87 : std_logic;
  signal gl_gr_lg_n_88, gl_gr_lg_n_89, gl_gr_lg_n_90, gl_gr_lg_n_91, gl_gr_lg_n_92 : std_logic;
  signal gl_gr_lg_n_93, gl_gr_lg_n_94, gl_gr_lg_n_95, gl_gr_lg_n_96, gl_gr_lg_n_97 : std_logic;
  signal gl_gr_lg_n_98, gl_gr_lg_n_99, gl_gr_lg_n_100, gl_gr_lg_n_101, gl_gr_lg_n_102 : std_logic;
  signal gl_gr_lg_n_103, gl_gr_lg_n_104, gl_gr_lg_n_105, gl_gr_lg_n_106, gl_gr_lg_n_107 : std_logic;
  signal gl_gr_lg_n_108, gl_gr_lg_n_109, gl_gr_lg_n_110, gl_gr_lg_n_111, gl_gr_lg_n_112 : std_logic;
  signal gl_gr_lg_n_113, gl_gr_lg_n_114, gl_gr_lg_n_115, gl_gr_lg_n_116, gl_gr_lg_n_117 : std_logic;
  signal gl_gr_lg_n_118, gl_gr_lg_n_155, gl_gr_lg_n_156, gl_ram_n_0, gl_ram_n_1 : std_logic;
  signal gl_ram_n_2, gl_ram_n_3, gl_ram_n_4, gl_ram_n_5, gl_ram_n_6 : std_logic;
  signal gl_ram_n_7, gl_ram_n_8, gl_ram_n_9, gl_ram_n_10, gl_ram_n_11 : std_logic;
  signal gl_ram_n_12, gl_ram_n_13, gl_ram_n_14, gl_ram_n_15, gl_ram_n_16 : std_logic;
  signal gl_ram_n_17, gl_ram_n_18, gl_ram_n_19, gl_ram_n_20, gl_ram_n_21 : std_logic;
  signal gl_ram_n_22, gl_ram_n_23, gl_ram_n_24, gl_ram_n_25, gl_ram_n_26 : std_logic;
  signal gl_ram_n_27, gl_ram_n_28, gl_ram_n_29, gl_ram_n_30, gl_ram_n_31 : std_logic;
  signal gl_ram_n_32, gl_ram_n_33, gl_ram_n_34, gl_ram_n_35, gl_ram_n_36 : std_logic;
  signal gl_ram_n_37, gl_ram_n_38, gl_ram_n_39, gl_ram_n_40, gl_ram_n_41 : std_logic;
  signal gl_ram_n_42, gl_ram_n_43, gl_ram_n_44, gl_ram_n_45, gl_ram_n_46 : std_logic;
  signal gl_ram_n_47, gl_ram_n_48, gl_ram_n_49, gl_ram_n_50, gl_ram_n_51 : std_logic;
  signal gl_ram_n_52, gl_ram_n_53, gl_ram_n_54, gl_ram_n_55, gl_ram_n_56 : std_logic;
  signal gl_ram_n_57, gl_ram_n_58, gl_ram_n_59, gl_ram_n_60, gl_ram_n_61 : std_logic;
  signal gl_ram_n_62, gl_ram_n_63, gl_ram_n_64, gl_ram_n_65, gl_ram_n_66 : std_logic;
  signal gl_ram_n_67, gl_ram_n_68, gl_ram_n_69, gl_ram_n_70, gl_ram_n_71 : std_logic;
  signal gl_ram_n_72, gl_ram_n_73, gl_ram_n_74, gl_ram_n_75, gl_ram_n_76 : std_logic;
  signal gl_ram_n_77, gl_ram_n_78, gl_ram_n_79, gl_ram_n_80, gl_ram_n_81 : std_logic;
  signal gl_ram_n_82, gl_ram_n_83, gl_ram_n_84, gl_ram_n_85, gl_ram_n_86 : std_logic;
  signal gl_ram_n_87, gl_ram_n_88, gl_ram_n_89, gl_ram_n_90, gl_ram_n_91 : std_logic;
  signal gl_ram_n_92, gl_ram_n_93, gl_ram_n_94, gl_ram_n_95, gl_ram_n_96 : std_logic;
  signal gl_ram_n_97, gl_ram_n_98, gl_ram_n_99, gl_ram_n_100, gl_ram_n_101 : std_logic;
  signal gl_ram_n_102, gl_ram_n_103, gl_ram_n_104, gl_ram_n_105, gl_ram_n_106 : std_logic;
  signal gl_ram_n_107, gl_ram_n_108, gl_ram_n_109, gl_ram_n_110, gl_ram_n_111 : std_logic;
  signal gl_ram_n_112, gl_ram_n_113, gl_ram_n_114, gl_ram_n_115, gl_ram_n_116 : std_logic;
  signal gl_ram_n_117, gl_ram_n_118, gl_ram_n_119, gl_ram_n_120, gl_ram_n_121 : std_logic;
  signal gl_ram_n_122, gl_ram_n_123, gl_ram_n_124, gl_ram_n_125, gl_ram_n_126 : std_logic;
  signal gl_ram_n_127, gl_ram_n_128, gl_ram_n_129, gl_ram_n_130, gl_ram_n_131 : std_logic;
  signal gl_ram_n_132, gl_ram_n_133, gl_ram_n_134, gl_ram_n_135, gl_ram_n_136 : std_logic;
  signal gl_ram_n_137, gl_ram_n_138, gl_ram_n_139, gl_ram_n_140, gl_ram_n_141 : std_logic;
  signal gl_ram_n_142, gl_ram_n_143, gl_ram_n_144, gl_ram_n_145, gl_ram_n_146 : std_logic;
  signal gl_ram_n_147, gl_ram_n_148, gl_ram_n_149, gl_ram_n_150, gl_ram_n_151 : std_logic;
  signal gl_ram_n_152, gl_ram_n_153, gl_ram_n_154, gl_ram_n_155, gl_ram_n_156 : std_logic;
  signal gl_ram_n_157, gl_ram_n_158, gl_ram_n_159, gl_ram_n_160, gl_ram_n_161 : std_logic;
  signal gl_ram_n_162, gl_ram_n_163, gl_ram_n_164, gl_ram_n_165, gl_ram_n_166 : std_logic;
  signal gl_ram_n_167, gl_ram_n_168, gl_ram_n_169, gl_ram_n_170, gl_ram_n_171 : std_logic;
  signal gl_ram_n_172, gl_ram_n_173, gl_ram_n_174, gl_ram_n_175, gl_ram_n_176 : std_logic;
  signal gl_ram_n_177, gl_ram_n_178, gl_ram_n_179, gl_ram_n_180, gl_ram_n_181 : std_logic;
  signal gl_ram_n_182, gl_ram_n_183, gl_ram_n_184, gl_ram_n_185, gl_ram_n_186 : std_logic;
  signal gl_ram_n_187, gl_ram_n_188, gl_ram_n_189, gl_ram_n_190, gl_ram_n_191 : std_logic;
  signal gl_ram_n_192, gl_ram_n_193, gl_ram_n_194, gl_ram_n_195, gl_ram_n_196 : std_logic;
  signal gl_ram_n_197, gl_ram_n_198, gl_ram_n_199, gl_ram_n_200, gl_ram_n_201 : std_logic;
  signal gl_ram_n_202, gl_ram_n_203, gl_ram_n_204, gl_ram_n_205, gl_ram_n_206 : std_logic;
  signal gl_ram_n_207, gl_ram_n_208, gl_ram_n_209, gl_ram_n_210, gl_ram_n_211 : std_logic;
  signal gl_ram_n_212, gl_ram_n_213, gl_ram_n_214, gl_ram_n_215, gl_ram_n_216 : std_logic;
  signal gl_ram_n_217, gl_ram_n_218, gl_ram_n_219, gl_ram_n_220, gl_ram_n_221 : std_logic;
  signal gl_ram_n_222, gl_ram_n_223, gl_ram_n_224, gl_ram_n_225, gl_ram_n_226 : std_logic;
  signal gl_ram_n_227, gl_ram_n_228, gl_ram_n_229, gl_ram_n_230, gl_ram_n_231 : std_logic;
  signal gl_ram_n_232, gl_ram_n_233, gl_ram_n_234, gl_ram_n_235, gl_ram_n_236 : std_logic;
  signal gl_ram_n_237, gl_ram_n_238, gl_ram_n_239, gl_ram_n_240, gl_ram_n_241 : std_logic;
  signal gl_ram_n_242, gl_ram_n_243, gl_ram_n_244, gl_ram_n_245, gl_ram_n_246 : std_logic;
  signal gl_ram_n_247, gl_ram_n_248, gl_ram_n_249, gl_ram_n_250, gl_ram_n_251 : std_logic;
  signal gl_ram_n_252, gl_ram_n_253, gl_ram_n_254, gl_ram_n_255, gl_ram_n_256 : std_logic;
  signal gl_ram_n_257, gl_ram_n_258, gl_ram_n_259, gl_ram_n_260, gl_ram_n_261 : std_logic;
  signal gl_ram_n_262, gl_ram_n_263, gl_ram_n_264, gl_ram_n_265, gl_ram_n_266 : std_logic;
  signal gl_ram_n_267, gl_ram_n_268, gl_ram_n_269, gl_ram_n_270, gl_ram_n_271 : std_logic;
  signal gl_ram_n_272, gl_ram_n_273, gl_ram_n_274, gl_ram_n_275, gl_ram_n_276 : std_logic;
  signal gl_ram_n_277, gl_ram_n_278, gl_ram_n_279, gl_ram_n_280, gl_ram_n_281 : std_logic;
  signal gl_ram_n_282, gl_ram_n_283, gl_ram_n_284, gl_ram_n_285, gl_ram_n_286 : std_logic;
  signal gl_ram_n_287, gl_ram_n_288, gl_ram_n_289, gl_ram_n_290, gl_ram_n_291 : std_logic;
  signal gl_ram_n_292, gl_ram_n_293, gl_ram_n_294, gl_ram_n_295, gl_ram_n_296 : std_logic;
  signal gl_ram_n_297, gl_ram_n_298, gl_ram_n_299, gl_ram_n_300, gl_ram_n_301 : std_logic;
  signal gl_ram_n_302, gl_ram_n_303, gl_ram_n_304, gl_ram_n_305, gl_ram_n_306 : std_logic;
  signal gl_ram_n_307, gl_ram_n_308, gl_ram_n_309, gl_ram_n_310, gl_ram_n_311 : std_logic;
  signal gl_ram_n_312, gl_ram_n_313, gl_ram_n_314, gl_ram_n_315, gl_ram_n_316 : std_logic;
  signal gl_ram_n_317, gl_ram_n_318, gl_ram_n_319, gl_ram_n_320, gl_ram_n_321 : std_logic;
  signal gl_ram_n_322, gl_ram_n_323, gl_ram_n_324, gl_ram_n_325, gl_ram_n_326 : std_logic;
  signal gl_ram_n_327, gl_ram_n_328, gl_ram_n_329, gl_ram_n_330, gl_ram_n_331 : std_logic;
  signal gl_ram_n_332, gl_ram_n_333, gl_ram_n_334, gl_ram_n_335, gl_ram_n_336 : std_logic;
  signal gl_ram_n_337, gl_ram_n_338, gl_ram_n_339, gl_ram_n_340, gl_ram_n_341 : std_logic;
  signal gl_ram_n_342, gl_ram_n_343, gl_ram_n_344, gl_ram_n_345, gl_ram_n_346 : std_logic;
  signal gl_ram_n_347, gl_ram_n_348, gl_ram_n_349, gl_ram_n_350, gl_ram_n_351 : std_logic;
  signal gl_ram_n_352, gl_ram_n_353, gl_ram_n_354, gl_ram_n_355, gl_ram_n_356 : std_logic;
  signal gl_ram_n_357, gl_ram_n_358, gl_ram_n_359, gl_ram_n_360, gl_ram_n_361 : std_logic;
  signal gl_ram_n_362, gl_ram_n_363, gl_ram_n_364, gl_ram_n_365, gl_ram_n_366 : std_logic;
  signal gl_ram_n_367, gl_ram_n_368, gl_ram_n_369, gl_ram_n_370, gl_ram_n_371 : std_logic;
  signal gl_ram_n_372, gl_ram_n_373, gl_ram_n_374, gl_ram_n_375, gl_ram_n_376 : std_logic;
  signal gl_ram_n_377, gl_ram_n_378, gl_ram_n_379, gl_ram_n_380, gl_ram_n_381 : std_logic;
  signal gl_ram_n_382, gl_ram_n_383, gl_ram_n_384, gl_ram_n_385, gl_ram_n_386 : std_logic;
  signal gl_ram_n_387, gl_ram_n_388, gl_ram_n_389, gl_ram_n_390, gl_ram_n_391 : std_logic;
  signal gl_ram_n_392, gl_ram_n_393, gl_ram_n_394, gl_ram_n_395, gl_ram_n_396 : std_logic;
  signal gl_ram_n_397, gl_ram_n_398, gl_ram_n_399, gl_ram_n_400, gl_ram_n_401 : std_logic;
  signal gl_ram_n_402, gl_ram_n_403, gl_ram_n_404, gl_ram_n_405, gl_ram_n_406 : std_logic;
  signal gl_ram_n_407, gl_ram_n_408, gl_ram_n_409, gl_ram_n_410, gl_ram_n_411 : std_logic;
  signal gl_ram_n_412, gl_ram_n_413, gl_ram_n_414, gl_ram_n_415, gl_ram_n_416 : std_logic;
  signal gl_ram_n_417, gl_ram_n_418, gl_ram_n_419, gl_ram_n_420, gl_ram_n_421 : std_logic;
  signal gl_ram_n_422, gl_ram_n_423, gl_ram_n_424, gl_ram_n_425, gl_ram_n_426 : std_logic;
  signal gl_ram_n_427, gl_ram_n_428, gl_ram_n_429, gl_ram_n_430, gl_ram_n_431 : std_logic;
  signal gl_ram_n_432, gl_ram_n_433, gl_ram_n_434, gl_ram_n_435, gl_ram_n_436 : std_logic;
  signal gl_ram_n_437, gl_ram_n_438, gl_ram_n_439, gl_ram_n_440, gl_ram_n_441 : std_logic;
  signal gl_ram_n_442, gl_ram_n_443, gl_ram_n_444, gl_ram_n_445, gl_ram_n_446 : std_logic;
  signal gl_ram_n_447, gl_ram_n_448, gl_ram_n_449, gl_ram_n_450, gl_ram_n_451 : std_logic;
  signal gl_ram_n_452, gl_ram_n_453, gl_ram_n_454, gl_ram_n_455, gl_ram_n_456 : std_logic;
  signal gl_ram_n_457, gl_ram_n_458, gl_ram_n_459, gl_ram_n_460, gl_ram_n_461 : std_logic;
  signal gl_ram_n_462, gl_ram_n_463, gl_ram_n_464, gl_ram_n_465, gl_ram_n_466 : std_logic;
  signal gl_ram_n_467, gl_ram_n_468, gl_ram_n_469, gl_ram_n_470, gl_ram_n_471 : std_logic;
  signal gl_ram_n_472, gl_ram_n_473, gl_ram_n_474, gl_ram_n_475, gl_ram_n_476 : std_logic;
  signal gl_ram_n_477, gl_ram_n_478, gl_ram_n_479, gl_ram_n_480, gl_ram_n_481 : std_logic;
  signal gl_ram_n_482, gl_ram_n_483, gl_ram_n_484, gl_ram_n_485, gl_ram_n_486 : std_logic;
  signal gl_ram_n_487, gl_ram_n_488, gl_ram_n_489, gl_ram_n_490, gl_ram_n_491 : std_logic;
  signal gl_ram_n_492, gl_ram_n_493, gl_ram_n_494, gl_ram_n_495, gl_ram_n_496 : std_logic;
  signal gl_ram_n_497, gl_ram_n_498, gl_ram_n_499, gl_ram_n_500, gl_ram_n_501 : std_logic;
  signal gl_ram_n_502, gl_ram_n_503, gl_ram_n_504, gl_ram_n_505, gl_ram_n_506 : std_logic;
  signal gl_ram_n_507, gl_ram_n_508, gl_ram_n_509, gl_ram_n_510, gl_ram_n_511 : std_logic;
  signal gl_ram_n_512, gl_ram_n_513, gl_ram_n_514, gl_ram_n_515, gl_ram_n_516 : std_logic;
  signal gl_ram_n_517, gl_ram_n_518, gl_ram_n_519, gl_ram_n_520, gl_ram_n_521 : std_logic;
  signal gl_ram_n_522, gl_ram_n_523, gl_ram_n_524, gl_ram_n_525, gl_ram_n_526 : std_logic;
  signal gl_ram_n_527, gl_ram_n_528, gl_ram_n_529, gl_ram_n_530, gl_ram_n_531 : std_logic;
  signal gl_ram_n_532, gl_ram_n_533, gl_ram_n_534, gl_ram_n_535, gl_ram_n_536 : std_logic;
  signal gl_ram_n_537, gl_ram_n_538, gl_ram_n_539, gl_ram_n_540, gl_ram_n_541 : std_logic;
  signal gl_ram_n_542, gl_ram_n_543, gl_ram_n_544, gl_ram_n_545, gl_ram_n_546 : std_logic;
  signal gl_ram_n_547, gl_ram_n_548, gl_ram_n_549, gl_ram_n_550, gl_ram_n_551 : std_logic;
  signal gl_ram_n_552, gl_ram_n_553, gl_ram_n_554, gl_ram_n_555, gl_ram_n_556 : std_logic;
  signal gl_ram_n_557, gl_ram_n_558, gl_ram_n_559, gl_ram_n_560, gl_ram_n_561 : std_logic;
  signal gl_ram_n_562, gl_ram_n_563, gl_ram_n_564, gl_ram_n_565, gl_ram_n_566 : std_logic;
  signal gl_ram_n_567, gl_ram_n_568, gl_ram_n_569, gl_ram_n_570, gl_ram_n_571 : std_logic;
  signal gl_ram_n_572, gl_ram_n_573, gl_ram_n_574, gl_ram_n_575, gl_ram_n_576 : std_logic;
  signal gl_ram_n_577, gl_ram_n_578, gl_ram_n_579, gl_ram_n_580, gl_ram_n_581 : std_logic;
  signal gl_ram_n_582, gl_ram_n_583, gl_ram_n_584, gl_ram_n_585, gl_ram_n_586 : std_logic;
  signal gl_ram_n_587, gl_ram_n_588, gl_ram_n_589, gl_ram_n_590, gl_ram_n_591 : std_logic;
  signal gl_ram_n_592, gl_ram_n_593, gl_ram_n_594, gl_ram_n_595, gl_ram_n_596 : std_logic;
  signal gl_ram_n_597, gl_ram_n_598, gl_ram_n_599, gl_ram_n_600, gl_ram_n_601 : std_logic;
  signal gl_ram_n_602, gl_ram_n_603, gl_ram_n_604, gl_ram_n_605, gl_ram_n_606 : std_logic;
  signal gl_ram_n_607, gl_ram_n_608, gl_ram_n_609, gl_ram_n_610, gl_ram_n_611 : std_logic;
  signal gl_ram_n_612, gl_ram_n_613, gl_ram_n_614, gl_ram_n_615, gl_ram_n_616 : std_logic;
  signal gl_ram_n_617, gl_ram_n_618, gl_ram_n_619, gl_ram_n_620, gl_ram_n_621 : std_logic;
  signal gl_ram_n_622, gl_ram_n_623, gl_ram_n_624, gl_ram_n_625, gl_ram_n_626 : std_logic;
  signal gl_ram_n_627, gl_ram_n_628, gl_ram_n_629, gl_ram_n_630, gl_ram_n_631 : std_logic;
  signal gl_ram_n_632, gl_ram_n_633, gl_ram_n_634, gl_ram_n_635, gl_ram_n_636 : std_logic;
  signal gl_ram_n_637, gl_ram_n_638, gl_ram_n_639, gl_ram_n_640, gl_ram_n_641 : std_logic;
  signal gl_ram_n_642, gl_ram_n_643, gl_ram_n_644, gl_ram_n_645, gl_ram_n_646 : std_logic;
  signal gl_ram_n_647, gl_ram_n_648, gl_ram_n_649, gl_ram_n_650, gl_ram_n_651 : std_logic;
  signal gl_ram_n_652, gl_ram_n_653, gl_ram_n_654, gl_ram_n_655, gl_ram_n_656 : std_logic;
  signal gl_ram_n_657, gl_ram_n_658, gl_ram_n_659, gl_ram_n_660, gl_ram_n_661 : std_logic;
  signal gl_ram_n_662, gl_ram_n_663, gl_ram_n_664, gl_ram_n_665, gl_ram_n_666 : std_logic;
  signal gl_ram_n_667, gl_ram_n_668, gl_ram_n_669, gl_ram_n_670, gl_ram_n_671 : std_logic;
  signal gl_ram_n_672, gl_ram_n_673, gl_ram_n_674, gl_ram_n_675, gl_ram_n_676 : std_logic;
  signal gl_ram_n_677, gl_ram_n_678, gl_ram_n_679, gl_ram_n_680, gl_ram_n_681 : std_logic;
  signal gl_ram_n_682, gl_ram_n_683, gl_ram_n_684, gl_ram_n_685, gl_ram_n_686 : std_logic;
  signal gl_ram_n_687, gl_ram_n_688, gl_ram_n_689, gl_ram_n_690, gl_ram_n_691 : std_logic;
  signal gl_ram_n_692, gl_ram_n_693, gl_ram_n_694, gl_ram_n_695, gl_ram_n_696 : std_logic;
  signal gl_ram_n_697, gl_ram_n_698, gl_ram_n_699, gl_ram_n_700, gl_ram_n_701 : std_logic;
  signal gl_ram_n_702, gl_ram_n_703, gl_ram_n_704, gl_ram_n_705, gl_ram_n_706 : std_logic;
  signal gl_ram_n_707, gl_ram_n_708, gl_ram_n_709, gl_ram_n_710, gl_ram_n_711 : std_logic;
  signal gl_ram_n_712, gl_ram_n_713, gl_ram_n_714, gl_ram_n_715, gl_ram_n_716 : std_logic;
  signal gl_ram_n_717, gl_ram_n_718, gl_ram_n_719, gl_ram_n_720, gl_ram_n_721 : std_logic;
  signal gl_ram_n_722, gl_ram_n_723, gl_ram_n_724, gl_ram_n_725, gl_ram_n_726 : std_logic;
  signal gl_ram_n_727, gl_ram_n_728, gl_ram_n_729, gl_ram_n_730, gl_ram_n_731 : std_logic;
  signal gl_ram_n_732, gl_ram_n_733, gl_ram_n_734, gl_ram_n_735, gl_ram_n_736 : std_logic;
  signal gl_ram_n_737, gl_ram_n_738, gl_ram_n_739, gl_ram_n_740, gl_ram_n_741 : std_logic;
  signal gl_ram_n_742, gl_ram_n_743, gl_ram_n_744, gl_ram_n_745, gl_ram_n_746 : std_logic;
  signal gl_ram_n_747, gl_ram_n_748, gl_ram_n_749, gl_ram_n_750, gl_ram_n_751 : std_logic;
  signal gl_ram_n_752, gl_ram_n_753, gl_ram_n_754, gl_ram_n_755, gl_ram_n_756 : std_logic;
  signal gl_ram_n_757, gl_ram_n_758, gl_ram_n_759, gl_ram_n_760, gl_ram_n_761 : std_logic;
  signal gl_ram_n_762, gl_ram_n_763, gl_ram_n_764, gl_ram_n_765, gl_ram_n_766 : std_logic;
  signal gl_ram_n_767, gl_ram_n_768, gl_ram_n_769, gl_ram_n_770, gl_ram_n_771 : std_logic;
  signal gl_ram_n_772, gl_ram_n_773, gl_ram_n_774, gl_ram_n_775, gl_ram_n_776 : std_logic;
  signal gl_ram_n_777, gl_ram_n_778, gl_ram_n_779, gl_ram_n_780, gl_ram_n_781 : std_logic;
  signal gl_ram_n_782, gl_ram_n_783, gl_ram_n_784, gl_ram_n_785, gl_ram_n_786 : std_logic;
  signal gl_ram_n_787, gl_ram_n_788, gl_ram_n_789, gl_ram_n_790, gl_ram_n_791 : std_logic;
  signal gl_ram_n_792, gl_ram_n_793, gl_ram_n_794, gl_ram_n_795, gl_ram_n_796 : std_logic;
  signal gl_ram_n_797, gl_ram_n_798, gl_ram_n_799, gl_ram_n_800, gl_ram_n_801 : std_logic;
  signal gl_ram_n_802, gl_ram_n_803, gl_ram_n_804, gl_ram_n_805, gl_ram_n_806 : std_logic;
  signal gl_ram_n_807, gl_ram_n_808, gl_ram_n_809, gl_ram_n_810, gl_ram_n_811 : std_logic;
  signal gl_ram_n_812, gl_ram_n_813, gl_ram_n_814, gl_ram_n_815, gl_ram_n_816 : std_logic;
  signal gl_ram_n_817, gl_ram_n_818, gl_ram_n_819, gl_ram_n_820, gl_ram_n_821 : std_logic;
  signal gl_ram_n_822, gl_ram_n_823, gl_ram_n_824, gl_ram_n_825, gl_ram_n_826 : std_logic;
  signal gl_ram_n_827, gl_ram_n_828, gl_ram_n_829, gl_ram_n_830, gl_ram_n_831 : std_logic;
  signal gl_ram_n_832, gl_ram_n_833, gl_ram_n_834, gl_ram_n_835, gl_ram_n_836 : std_logic;
  signal gl_ram_n_837, gl_ram_n_838, gl_ram_n_839, gl_ram_n_840, gl_ram_n_841 : std_logic;
  signal gl_ram_n_842, gl_ram_n_843, gl_ram_n_844, gl_ram_n_845, gl_ram_n_846 : std_logic;
  signal gl_ram_n_847, gl_ram_n_848, gl_ram_n_849, gl_ram_n_850, gl_ram_n_851 : std_logic;
  signal gl_ram_n_852, gl_ram_n_853, gl_ram_n_854, gl_ram_n_855, gl_ram_n_856 : std_logic;
  signal gl_ram_n_857, gl_ram_n_858, gl_ram_n_859, gl_ram_n_860, gl_ram_n_861 : std_logic;
  signal gl_ram_n_862, gl_ram_n_863, gl_ram_n_864, gl_ram_n_865, gl_ram_n_866 : std_logic;
  signal gl_ram_n_867, gl_ram_n_868, gl_ram_n_869, gl_ram_n_870, gl_ram_n_871 : std_logic;
  signal gl_ram_n_872, gl_ram_n_873, gl_ram_n_874, gl_ram_n_875, gl_ram_n_876 : std_logic;
  signal gl_ram_n_877, gl_ram_n_878, gl_ram_n_879, gl_ram_n_880, gl_ram_n_881 : std_logic;
  signal gl_ram_n_882, gl_ram_n_883, gl_ram_n_884, gl_ram_n_885, gl_ram_n_886 : std_logic;
  signal gl_ram_n_887, gl_ram_n_888, gl_ram_n_889, gl_ram_n_890, gl_ram_n_891 : std_logic;
  signal gl_ram_n_892, gl_ram_n_893, gl_ram_n_894, gl_ram_n_895, gl_ram_n_896 : std_logic;
  signal gl_ram_n_897, gl_ram_n_898, gl_ram_n_899, gl_ram_n_900, gl_ram_n_901 : std_logic;
  signal gl_ram_n_902, gl_ram_n_903, gl_ram_n_904, gl_ram_n_905, gl_ram_n_906 : std_logic;
  signal gl_ram_n_907, gl_ram_n_908, gl_ram_n_909, gl_ram_n_910, gl_ram_n_911 : std_logic;
  signal gl_ram_n_912, gl_ram_n_913, gl_ram_n_914, gl_ram_n_915, gl_ram_n_916 : std_logic;
  signal gl_ram_n_917, gl_ram_n_918, gl_ram_n_919, gl_ram_n_920, gl_ram_n_921 : std_logic;
  signal gl_ram_n_922, gl_ram_n_923, gl_ram_n_924, gl_ram_n_925, gl_ram_n_926 : std_logic;
  signal gl_ram_n_927, gl_ram_n_928, gl_ram_n_929, gl_ram_n_930, gl_ram_n_931 : std_logic;
  signal gl_ram_n_932, gl_ram_n_933, gl_ram_n_934, gl_ram_n_935, gl_ram_n_936 : std_logic;
  signal gl_ram_n_937, gl_ram_n_938, gl_ram_n_939, gl_ram_n_940, gl_ram_n_941 : std_logic;
  signal gl_ram_n_942, gl_ram_n_943, gl_ram_n_944, gl_ram_n_945, gl_ram_n_946 : std_logic;
  signal gl_ram_n_947, gl_ram_n_948, gl_ram_n_949, gl_ram_n_950, gl_ram_n_951 : std_logic;
  signal gl_ram_n_952, gl_ram_n_953, gl_ram_n_954, gl_ram_n_955, gl_ram_n_956 : std_logic;
  signal gl_ram_n_957, gl_ram_n_958, gl_ram_n_959, gl_ram_n_960, gl_ram_n_961 : std_logic;
  signal gl_ram_n_962, gl_ram_n_963, gl_ram_n_964, gl_ram_n_965, gl_ram_n_966 : std_logic;
  signal gl_ram_n_967, gl_ram_n_968, gl_ram_n_969, gl_ram_n_970, gl_ram_n_971 : std_logic;
  signal gl_ram_n_972, gl_ram_n_973, gl_ram_n_974, gl_ram_n_975, gl_ram_n_976 : std_logic;
  signal gl_ram_n_977, gl_ram_n_978, gl_ram_n_979, gl_ram_n_980, gl_ram_n_981 : std_logic;
  signal gl_ram_n_982, gl_ram_n_983, gl_ram_n_984, gl_ram_n_985, gl_ram_n_986 : std_logic;
  signal gl_ram_n_987, gl_ram_n_988, gl_ram_n_989, gl_ram_n_990, gl_ram_n_991 : std_logic;
  signal gl_ram_n_992, gl_ram_n_993, gl_ram_n_994, gl_ram_n_995, gl_ram_n_996 : std_logic;
  signal gl_ram_n_997, gl_ram_n_998, gl_ram_n_999, gl_ram_n_1000, gl_ram_n_1001 : std_logic;
  signal gl_ram_n_1002, gl_ram_n_1003, gl_ram_n_1004, gl_ram_n_1005, gl_ram_n_1006 : std_logic;
  signal gl_ram_n_1007, gl_ram_n_1008, gl_ram_n_1009, gl_ram_n_1010, gl_ram_n_1011 : std_logic;
  signal gl_ram_n_1012, gl_ram_n_1013, gl_ram_n_1014, gl_ram_n_1015, gl_ram_n_1016 : std_logic;
  signal gl_ram_n_1017, gl_ram_n_1018, gl_ram_n_1019, gl_ram_n_1020, gl_ram_n_1021 : std_logic;
  signal gl_ram_n_1022, gl_ram_n_1023, gl_ram_n_1024, gl_ram_n_1025, gl_ram_n_1026 : std_logic;
  signal gl_ram_n_1027, gl_ram_n_1028, gl_ram_n_1029, gl_ram_n_1030, gl_ram_n_1031 : std_logic;
  signal gl_ram_n_1032, gl_ram_n_1033, gl_ram_n_1034, gl_ram_n_1035, gl_ram_n_1036 : std_logic;
  signal gl_ram_n_1037, gl_ram_n_1038, gl_ram_n_1039, gl_ram_n_1040, gl_ram_n_1041 : std_logic;
  signal gl_ram_n_1042, gl_ram_n_1043, gl_ram_n_1044, gl_ram_n_1045, gl_ram_n_1046 : std_logic;
  signal gl_ram_n_1047, gl_ram_n_1048, gl_ram_n_1049, gl_ram_n_1050, gl_ram_n_1051 : std_logic;
  signal gl_ram_n_1052, gl_ram_n_1053, gl_ram_n_1054, gl_ram_n_1055, gl_ram_n_1056 : std_logic;
  signal gl_ram_n_1057, gl_ram_n_1058, gl_ram_n_1059, gl_rom_n_0, gl_rom_n_1 : std_logic;
  signal gl_rom_n_2, gl_rom_n_3, gl_rom_n_4, gl_rom_n_5, gl_rom_n_6 : std_logic;
  signal gl_rom_n_7, gl_rom_n_8, gl_rom_n_9, gl_rom_n_10, gl_rom_n_11 : std_logic;
  signal gl_rom_n_12, gl_rom_n_13, gl_rom_n_14, gl_rom_n_15, gl_rom_n_16 : std_logic;
  signal gl_rom_n_17, gl_rom_n_18, gl_rom_n_19, gl_rom_n_20, gl_rom_n_21 : std_logic;
  signal gl_rom_n_22, gl_rom_n_23, gl_rom_n_24, gl_rom_n_25, gl_rom_n_26 : std_logic;
  signal gl_rom_n_27, gl_rom_n_28, gl_rom_n_29, gl_rom_n_30, gl_rom_n_31 : std_logic;
  signal gl_rom_n_32, gl_rom_n_33, gl_rom_n_34, gl_rom_n_35, gl_rom_n_36 : std_logic;
  signal gl_rom_n_37, gl_rom_n_38, gl_rom_n_39, gl_rom_n_40, gl_rom_n_41 : std_logic;
  signal gl_rom_n_42, gl_rom_n_43, gl_rom_n_44, gl_rom_n_45, gl_rom_n_46 : std_logic;
  signal gl_rom_n_47, gl_rom_n_48, gl_rom_n_49, gl_rom_n_50, gl_rom_n_51 : std_logic;
  signal gl_rom_n_52, gl_rom_n_53, gl_rom_n_54, gl_rom_n_55, gl_rom_n_56 : std_logic;
  signal gl_rom_n_57, gl_rom_n_58, gl_rom_n_59, gl_rom_n_60, gl_rom_n_61 : std_logic;
  signal gl_rom_n_62, gl_rom_n_63, gl_rom_n_64, gl_rom_n_65, gl_rom_n_66 : std_logic;
  signal gl_rom_n_67, gl_rom_n_68, gl_rom_n_69, gl_rom_n_70, gl_rom_n_71 : std_logic;
  signal gl_rom_n_72, gl_rom_n_73, gl_rom_n_74, gl_rom_n_75, gl_rom_n_76 : std_logic;
  signal gl_rom_n_77, gl_rom_n_78, gl_rom_n_79, gl_rom_n_80, gl_rom_n_81 : std_logic;
  signal gl_rom_n_82, gl_rom_n_83, gl_rom_n_84, gl_rom_n_85, gl_rom_n_86 : std_logic;
  signal gl_rom_n_87, gl_rom_n_88, gl_rom_n_89, gl_rom_n_90, gl_rom_n_91 : std_logic;
  signal gl_rom_n_92, gl_rom_n_93, gl_rom_n_94, gl_rom_n_95, gl_rom_n_96 : std_logic;
  signal gl_rom_n_97, gl_rom_n_98, gl_rom_n_99, gl_rom_n_100, gl_rom_n_101 : std_logic;
  signal gl_rom_n_102, gl_rom_n_103, gl_rom_n_104, gl_rom_n_105, gl_rom_n_106 : std_logic;
  signal gl_rom_n_107, gl_rom_n_108, gl_rom_n_109, gl_rom_n_110, gl_rom_n_111 : std_logic;
  signal gl_rom_n_112, gl_rom_n_113, gl_rom_n_114, gl_rom_n_115, gl_rom_n_116 : std_logic;
  signal gl_rom_n_117, gl_rom_n_118, gl_rom_n_119, gl_rom_n_120, gl_rom_n_121 : std_logic;
  signal gl_rom_n_122, gl_rom_n_123, gl_rom_n_124, gl_rom_n_125, gl_rom_n_126 : std_logic;
  signal gl_rom_n_127, gl_rom_n_128, gl_rom_n_129, gl_rom_n_130, gl_rom_n_131 : std_logic;
  signal gl_rom_n_132, gl_rom_n_133, gl_rom_n_134, gl_rom_n_135, gl_rom_n_136 : std_logic;
  signal gl_rom_n_137, gl_rom_n_138, gl_rom_n_139, gl_rom_n_140, gl_rom_n_141 : std_logic;
  signal gl_rom_n_142, gl_rom_n_143, gl_rom_n_144, gl_rom_n_145, gl_rom_n_146 : std_logic;
  signal gl_rom_n_147, gl_rom_n_148, gl_rom_n_149, gl_rom_n_150, gl_rom_n_151 : std_logic;
  signal gl_rom_n_152, gl_rom_n_153, gl_rom_n_154, gl_rom_n_155, gl_rom_n_156 : std_logic;
  signal gl_rom_n_157, gl_rom_n_158, gl_rom_n_159, gl_rom_n_160, gl_rom_n_161 : std_logic;
  signal gl_rom_n_162, gl_rom_n_163, gl_rom_n_164, gl_rom_n_165, gl_rom_n_166 : std_logic;
  signal gl_rom_n_167, gl_rom_n_168, gl_rom_n_169, gl_rom_n_170, gl_rom_n_171 : std_logic;
  signal gl_rom_n_172, gl_rom_n_173, gl_rom_n_174, gl_rom_n_175, gl_rom_n_176 : std_logic;
  signal gl_rom_n_177, gl_rom_n_178, gl_rom_n_179, gl_rom_n_180, gl_rom_n_181 : std_logic;
  signal gl_rom_n_182, gl_rom_n_183, gl_rom_n_184, gl_rom_n_185, gl_rom_n_186 : std_logic;
  signal gl_rom_n_187, gl_rom_n_188, gl_rom_n_189, gl_rom_n_190, gl_rom_n_191 : std_logic;
  signal gl_rom_n_192, gl_rom_n_193, gl_rom_n_194, gl_rom_n_195, gl_rom_n_196 : std_logic;
  signal gl_rom_n_197, gl_rom_n_198, gl_rom_n_199, gl_rom_n_200, gl_rom_n_201 : std_logic;
  signal gl_rom_n_202, gl_rom_n_203, gl_rom_n_204, gl_rom_n_205, gl_rom_n_206 : std_logic;
  signal gl_rom_n_207, gl_rom_n_208, gl_rom_n_209, gl_rom_n_210, gl_rom_n_211 : std_logic;
  signal gl_rom_n_212, gl_rom_n_213, gl_rom_n_214, gl_rom_n_215, gl_rom_n_216 : std_logic;
  signal gl_rom_n_217, gl_rom_n_218, gl_rom_n_219, gl_rom_n_220, gl_rom_n_221 : std_logic;
  signal gl_rom_n_222, gl_rom_n_223, gl_rom_n_224, gl_rom_n_225, gl_rom_n_226 : std_logic;
  signal gl_rom_n_227, gl_rom_n_228, gl_rom_n_229, gl_rom_n_230, gl_rom_n_231 : std_logic;
  signal gl_rom_n_232, gl_rom_n_233, gl_rom_n_234, gl_rom_n_235, gl_rom_n_236 : std_logic;
  signal gl_rom_n_237, gl_rom_n_238, gl_rom_n_239, gl_rom_n_240, gl_rom_n_241 : std_logic;
  signal gl_rom_n_242, gl_rom_n_243, gl_rom_n_244, gl_rom_n_245, gl_rom_n_246 : std_logic;
  signal gl_rom_n_247, gl_rom_n_248, gl_rom_n_249, gl_rom_n_250, gl_rom_n_251 : std_logic;
  signal gl_rom_n_252, gl_rom_n_253, gl_rom_n_254, gl_rom_n_255, gl_rom_n_256 : std_logic;
  signal gl_rom_n_257, gl_rom_n_258, gl_rom_n_259, gl_rom_n_260, gl_rom_n_261 : std_logic;
  signal gl_rom_n_262, gl_rom_n_263, gl_rom_n_264, gl_rom_n_265, gl_rom_n_266 : std_logic;
  signal gl_rom_n_267, gl_rom_n_268, gl_rom_n_269, gl_rom_n_270, gl_rom_n_271 : std_logic;
  signal gl_rom_n_272, gl_rom_n_273, gl_rom_n_274, gl_rom_n_275, gl_rom_n_276 : std_logic;
  signal gl_rom_n_277, gl_rom_n_278, gl_rom_n_279, gl_rom_n_280, gl_rom_n_281 : std_logic;
  signal gl_rom_n_282, gl_rom_n_283, gl_rom_n_284, gl_rom_n_285, gl_rom_n_286 : std_logic;
  signal gl_rom_n_287, gl_rom_n_288, gl_rom_n_289, gl_rom_n_290, gl_rom_n_291 : std_logic;
  signal gl_rom_n_292, gl_rom_n_293, gl_rom_n_294, gl_rom_n_295, gl_rom_n_296 : std_logic;
  signal gl_rom_n_297, gl_rom_n_298, gl_rom_n_299, gl_rom_n_300, gl_rom_n_301 : std_logic;
  signal gl_rom_n_302, gl_rom_n_303, gl_rom_n_304, gl_rom_n_305, gl_rom_n_306 : std_logic;
  signal gl_rom_n_307, gl_rom_n_308, gl_rom_n_309, gl_rom_n_310, gl_rom_n_311 : std_logic;
  signal gl_rom_n_312, gl_rom_n_313, gl_rom_n_314, gl_rom_n_315, gl_rom_n_316 : std_logic;
  signal gl_rom_n_317, gl_rom_n_318, gl_rom_n_319, gl_rom_n_320, gl_rom_n_321 : std_logic;
  signal gl_rom_n_322, gl_rom_n_323, gl_rom_n_324, gl_rom_n_325, gl_rom_n_326 : std_logic;
  signal gl_rom_n_327, gl_rom_n_328, gl_rom_n_329, gl_rom_n_330, gl_rom_n_331 : std_logic;
  signal gl_rom_n_332, gl_rom_n_333, gl_rom_n_334, gl_rom_n_335, gl_rom_n_336 : std_logic;
  signal gl_rom_n_337, gl_rom_n_338, gl_rom_n_339, gl_rom_n_340, gl_rom_n_341 : std_logic;
  signal gl_rom_n_342, gl_rom_n_343, gl_rom_n_344, gl_rom_n_345, gl_rom_n_346 : std_logic;
  signal gl_rom_n_347, gl_rom_n_348, gl_rom_n_349, gl_rom_n_350, gl_rom_n_351 : std_logic;
  signal gl_rom_n_352, gl_rom_n_353, gl_rom_n_354, gl_rom_n_355, gl_rom_n_356 : std_logic;
  signal gl_rom_n_357, gl_rom_n_358, gl_rom_n_359, gl_rom_n_360, gl_rom_n_361 : std_logic;
  signal gl_rom_n_362, gl_rom_n_363, gl_rom_n_364, gl_rom_n_365, gl_rom_n_366 : std_logic;
  signal gl_rom_n_367, gl_rom_n_368, gl_rom_n_369, gl_rom_n_370, gl_rom_n_371 : std_logic;
  signal gl_rom_n_372, gl_rom_n_373, gl_rom_n_374, gl_rom_n_375, gl_rom_n_376 : std_logic;
  signal gl_rom_n_377, gl_rom_n_378, gl_rom_n_379, gl_rom_n_380, gl_rom_n_381 : std_logic;
  signal gl_rom_n_382, gl_rom_n_383, gl_rom_n_384, gl_rom_n_385, gl_rom_n_386 : std_logic;
  signal gl_rom_n_387, gl_rom_n_388, gl_rom_n_389, gl_rom_n_390, gl_rom_n_391 : std_logic;
  signal gl_rom_n_392, gl_rom_n_393, gl_rom_n_394, gl_rom_n_395, gl_rom_n_396 : std_logic;
  signal gl_rom_n_397, gl_rom_n_398, gl_rom_n_399, gl_rom_n_400, gl_rom_n_401 : std_logic;
  signal gl_rom_n_402, gl_rom_n_403, gl_rom_n_404, gl_rom_n_405, gl_rom_n_406 : std_logic;
  signal gl_rom_n_407, gl_rom_n_408, gl_rom_n_409, gl_rom_n_410, gl_rom_n_411 : std_logic;
  signal gl_rom_n_412, gl_rom_n_413, gl_rom_n_414, gl_rom_n_415, gl_rom_n_416 : std_logic;
  signal gl_rom_n_417, gl_rom_n_418, gl_rom_n_419, gl_rom_n_420, gl_rom_n_421 : std_logic;
  signal gl_rom_n_422, gl_rom_n_423, gl_rom_n_424, gl_rom_n_425, gl_rom_n_426 : std_logic;
  signal gl_rom_n_427, gl_rom_n_428, gl_rom_n_429, gl_rom_n_430, gl_rom_n_431 : std_logic;
  signal gl_rom_n_432, gl_rom_n_433, gl_rom_n_434, gl_rom_n_435, gl_rom_n_436 : std_logic;
  signal gl_rom_n_437, gl_rom_n_438, gl_rom_n_439, gl_rom_n_440, gl_rom_n_441 : std_logic;
  signal gl_rom_n_442, gl_rom_n_443, gl_rom_n_444, gl_rom_n_445, gl_rom_n_446 : std_logic;
  signal gl_rom_n_447, gl_rom_n_448, gl_rom_n_449, gl_rom_n_450, gl_rom_n_451 : std_logic;
  signal gl_rom_n_452, gl_rom_n_453, gl_rom_n_454, gl_rom_n_455, gl_rom_n_456 : std_logic;
  signal gl_rom_n_457, gl_rom_n_458, gl_rom_n_459, gl_rom_n_460, gl_rom_n_461 : std_logic;
  signal gl_rom_n_462, gl_rom_n_463, gl_rom_n_464, gl_rom_n_465, gl_rom_n_466 : std_logic;
  signal gl_rom_n_467, gl_rom_n_468, gl_rom_n_469, gl_rom_n_470, gl_rom_n_471 : std_logic;
  signal gl_rom_n_472, gl_rom_n_473, gl_rom_n_474, gl_rom_n_475, gl_rom_n_476 : std_logic;
  signal gl_rom_n_477, gl_rom_n_478, gl_rom_n_479, gl_rom_n_480, gl_rom_n_481 : std_logic;
  signal gl_rom_n_482, gl_rom_n_483, gl_rom_n_484, gl_rom_n_485, gl_rom_n_486 : std_logic;
  signal gl_rom_n_487, gl_rom_n_488, gl_rom_n_489, gl_rom_n_490, gl_rom_n_491 : std_logic;
  signal gl_rom_n_492, gl_rom_n_493, gl_rom_n_494, gl_rom_n_495, gl_rom_n_496 : std_logic;
  signal gl_rom_n_497, gl_rom_n_498, gl_rom_n_499, gl_rom_n_500, gl_rom_n_501 : std_logic;
  signal gl_rom_n_502, gl_rom_n_503, gl_rom_n_504, gl_rom_n_505, gl_rom_n_506 : std_logic;
  signal gl_rom_n_507, gl_rom_n_508, gl_rom_n_509, gl_rom_n_510, gl_rom_n_511 : std_logic;
  signal gl_rom_n_512, gl_rom_n_513, gl_rom_n_514, gl_rom_n_515, gl_rom_n_516 : std_logic;
  signal gl_rom_n_517, gl_rom_n_518, gl_rom_n_519, gl_rom_n_520, gl_rom_n_521 : std_logic;
  signal gl_rom_n_522, gl_rom_n_523, gl_rom_n_524, gl_rom_n_525, gl_rom_n_526 : std_logic;
  signal gl_rom_n_527, gl_rom_n_528, gl_rom_n_529, gl_rom_n_530, gl_rom_n_531 : std_logic;
  signal gl_rom_n_532, gl_rom_n_533, gl_rom_n_534, gl_rom_n_535, gl_rom_n_536 : std_logic;
  signal gl_rom_n_537, gl_rom_n_538, gl_rom_n_539, gl_rom_n_540, gl_rom_n_541 : std_logic;
  signal gl_rom_n_542, gl_rom_n_543, gl_rom_n_544, gl_rom_n_545, gl_rom_n_546 : std_logic;
  signal gl_rom_n_547, gl_rom_n_548, gl_rom_n_549, gl_rom_n_550, gl_rom_n_551 : std_logic;
  signal gl_rom_n_552, gl_rom_n_553, gl_rom_n_554, gl_rom_n_555, gl_rom_n_556 : std_logic;
  signal gl_rom_n_557, gl_rom_n_558, gl_rom_n_559, gl_rom_n_560, gl_rom_n_561 : std_logic;
  signal gl_rom_n_562, gl_rom_n_563, gl_rom_n_564, gl_rom_n_565, gl_rom_n_566 : std_logic;
  signal gl_rom_n_567, gl_rom_n_568, gl_rom_n_569, gl_rom_n_570, gl_rom_n_571 : std_logic;
  signal gl_rom_n_572, gl_rom_n_573, gl_rom_n_574, gl_rom_n_575, gl_rom_n_576 : std_logic;
  signal gl_rom_n_577, gl_rom_n_578, gl_rom_n_579, gl_rom_n_580, gl_rom_n_581 : std_logic;
  signal gl_rom_n_582, gl_rom_n_583, gl_rom_n_584, gl_rom_n_585, gl_rom_n_586 : std_logic;
  signal gl_rom_n_587, gl_rom_n_588, gl_rom_n_589, gl_rom_n_590, gl_rom_n_591 : std_logic;
  signal gl_rom_n_592, gl_rom_n_593, gl_rom_n_594, gl_rom_n_595, gl_rom_n_596 : std_logic;
  signal gl_rom_n_597, gl_rom_n_598, gl_rom_n_599, gl_rom_n_600, gl_rom_n_601 : std_logic;
  signal gl_rom_n_602, gl_rom_n_603, gl_rom_n_604, gl_rom_n_605, gl_rom_n_606 : std_logic;
  signal gl_rom_n_607, gl_rom_n_608, gl_rom_n_609, gl_rom_n_610, gl_rom_n_611 : std_logic;
  signal gl_rom_n_612, gl_rom_n_613, gl_rom_n_614, gl_rom_n_615, gl_rom_n_616 : std_logic;
  signal gl_rom_n_617, gl_rom_n_618, gl_rom_n_619, gl_rom_n_620, gl_rom_n_621 : std_logic;
  signal gl_rom_n_622, gl_rom_n_623, gl_rom_n_624, gl_rom_n_625, gl_rom_n_626 : std_logic;
  signal gl_rom_n_627, gl_rom_n_628, gl_rom_n_629, gl_rom_n_630, gl_rom_n_631 : std_logic;
  signal gl_rom_n_632, gl_rom_n_633, gl_rom_n_634, gl_rom_n_635, gl_rom_n_636 : std_logic;
  signal gl_rom_n_637, gl_rom_n_638, gl_rom_n_639, gl_rom_n_640, gl_rom_n_641 : std_logic;
  signal gl_rom_n_642, gl_rom_n_643, gl_rom_n_644, gl_rom_n_645, gl_rom_n_646 : std_logic;
  signal gl_rom_n_647, gl_rom_n_648, gl_rom_n_649, gl_rom_n_650, gl_rom_n_651 : std_logic;
  signal gl_rom_n_652, gl_rom_n_653, gl_rom_n_654, gl_rom_n_655, gl_rom_n_656 : std_logic;
  signal gl_rom_n_657, gl_rom_n_658, gl_rom_n_659, gl_rom_n_660, gl_rom_n_661 : std_logic;
  signal gl_rom_n_662, gl_rom_n_663, gl_rom_n_664, gl_rom_n_665, gl_rom_n_666 : std_logic;
  signal gl_rom_n_667, gl_rom_n_668, gl_rom_n_669, gl_rom_n_670, gl_rom_n_671 : std_logic;
  signal gl_rom_n_672, gl_rom_n_673, gl_rom_n_674, gl_rom_n_675, gl_rom_n_676 : std_logic;
  signal gl_rom_n_677, gl_rom_n_678, gl_rom_n_679, gl_rom_n_680, gl_rom_n_681 : std_logic;
  signal gl_rom_n_682, gl_rom_n_683, gl_rom_n_684, gl_rom_n_685, gl_rom_n_686 : std_logic;
  signal gl_rom_n_687, gl_rom_n_688, gl_rom_n_689, gl_rom_n_690, gl_rom_n_691 : std_logic;
  signal gl_rom_n_692, gl_rom_n_693, gl_rom_n_694, gl_rom_n_695, gl_rom_n_696 : std_logic;
  signal gl_rom_n_697, gl_rom_n_698, gl_rom_n_699, gl_rom_n_700, gl_rom_n_701 : std_logic;
  signal gl_rom_n_702, gl_rom_n_703, gl_rom_n_704, gl_rom_n_705, gl_rom_n_706 : std_logic;
  signal gl_rom_n_707, gl_rom_n_708, gl_rom_n_709, gl_rom_n_710, gl_rom_n_711 : std_logic;
  signal gl_rom_n_712, gl_rom_n_713, gl_rom_n_714, gl_rom_n_715, gl_rom_n_716 : std_logic;
  signal gl_rom_n_717, gl_rom_n_718, gl_rom_n_719, gl_rom_n_720, gl_rom_n_721 : std_logic;
  signal gl_rom_n_722, gl_rom_n_723, gl_rom_n_724, gl_rom_n_725, gl_rom_n_726 : std_logic;
  signal gl_rom_n_727, gl_rom_n_728, gl_rom_n_729, gl_rom_n_730, gl_rom_n_731 : std_logic;
  signal gl_rom_n_732, gl_rom_n_733, gl_rom_n_734, gl_rom_n_735, gl_rom_n_736 : std_logic;
  signal gl_rom_n_737, gl_rom_n_738, gl_rom_n_739, gl_rom_n_740, gl_rom_n_741 : std_logic;
  signal gl_rom_n_742, gl_rom_n_743, gl_rom_n_744, gl_rom_n_745, gl_rom_n_746 : std_logic;
  signal gl_rom_n_747, gl_rom_n_748, gl_rom_n_749, gl_rom_n_750, gl_rom_n_751 : std_logic;
  signal gl_rom_n_752, gl_rom_n_753, gl_rom_n_754, gl_rom_n_755, gl_rom_n_756 : std_logic;
  signal gl_rom_n_757, gl_rom_n_758, gl_rom_n_759, gl_rom_n_760, gl_rom_n_761 : std_logic;
  signal gl_rom_n_762, gl_rom_n_763, gl_rom_n_764, gl_rom_n_765, gl_rom_n_766 : std_logic;
  signal gl_rom_n_767, gl_rom_n_768, gl_rom_n_769, gl_rom_n_770, gl_rom_n_771 : std_logic;
  signal gl_rom_n_772, gl_rom_n_773, gl_rom_n_774, gl_rom_n_775, gl_rom_n_776 : std_logic;
  signal gl_rom_n_777, gl_rom_n_778, gl_rom_n_779, gl_rom_n_780, gl_rom_n_781 : std_logic;
  signal gl_rom_n_782, gl_rom_n_783, gl_rom_n_784, gl_rom_n_785, gl_rom_n_786 : std_logic;
  signal gl_rom_n_787, gl_rom_n_788, gl_rom_n_789, gl_rom_n_790, gl_rom_n_791 : std_logic;
  signal gl_rom_n_792, gl_rom_n_793, gl_rom_n_794, gl_rom_n_795, gl_rom_n_796 : std_logic;
  signal gl_rom_n_797, gl_rom_n_798, gl_rom_n_799, gl_rom_n_800, gl_rom_n_801 : std_logic;
  signal gl_rom_n_802, gl_rom_n_803, gl_rom_n_804, gl_rom_n_805, gl_rom_n_806 : std_logic;
  signal gl_rom_n_807, gl_rom_n_808, gl_rom_n_809, gl_rom_n_810, gl_rom_n_811 : std_logic;
  signal gl_rom_n_812, gl_rom_n_813, gl_rom_n_814, gl_rom_n_815, gl_rom_n_816 : std_logic;
  signal gl_rom_n_817, gl_rom_n_818, gl_rom_n_819, gl_rom_n_820, gl_rom_n_821 : std_logic;
  signal gl_rom_n_822, gl_rom_n_823, gl_rom_n_824, gl_rom_n_825, gl_rom_n_826 : std_logic;
  signal gl_rom_n_827, gl_rom_n_828, gl_rom_n_829, gl_rom_n_830, gl_rom_n_831 : std_logic;
  signal gl_rom_n_832, gl_rom_n_833, gl_rom_n_834, gl_rom_n_835, gl_rom_n_836 : std_logic;
  signal gl_rom_n_837, gl_rom_n_838, gl_rom_n_839, gl_rom_n_840, gl_rom_n_841 : std_logic;
  signal gl_rom_n_842, gl_rom_n_843, gl_rom_n_844, gl_rom_n_845, gl_rom_n_846 : std_logic;
  signal gl_rom_n_847, gl_rom_n_848, gl_rom_n_849, gl_rom_n_850, gl_rom_n_851 : std_logic;
  signal gl_rom_n_852, gl_rom_n_853, gl_rom_n_854, gl_rom_n_855, gl_rom_n_856 : std_logic;
  signal gl_rom_n_857, gl_rom_n_858, gl_rom_n_859, gl_rom_n_860, gl_rom_n_861 : std_logic;
  signal gl_rom_n_862, gl_rom_n_863, gl_rom_n_864, gl_rom_n_865, gl_rom_n_866 : std_logic;
  signal gl_rom_n_867, gl_rom_n_868, gl_rom_n_869, gl_rom_n_870, gl_rom_n_871 : std_logic;
  signal gl_rom_n_872, gl_rom_n_873, gl_rom_n_874, gl_rom_n_875, gl_rom_n_876 : std_logic;
  signal gl_rom_n_877, gl_rom_n_878, gl_rom_n_879, gl_rom_n_880, gl_rom_n_881 : std_logic;
  signal gl_rom_n_882, gl_rom_n_883, gl_rom_n_884, gl_rom_n_885, gl_rom_n_886 : std_logic;
  signal gl_rom_n_887, gl_rom_n_888, gl_rom_n_889, gl_rom_n_890, gl_rom_n_891 : std_logic;
  signal gl_rom_n_892, gl_rom_n_893, gl_rom_n_894, gl_rom_n_895, gl_rom_n_896 : std_logic;
  signal gl_rom_n_897, gl_rom_n_898, gl_rom_n_899, gl_rom_n_900, gl_rom_n_901 : std_logic;
  signal gl_rom_n_902, gl_rom_n_903, gl_rom_n_904, gl_rom_n_905, gl_rom_n_906 : std_logic;
  signal gl_rom_n_907, gl_rom_n_908, gl_rom_n_909, gl_rom_n_910, gl_rom_n_911 : std_logic;
  signal gl_rom_n_912, gl_rom_n_913, gl_rom_n_914, gl_rom_n_915, gl_rom_n_916 : std_logic;
  signal gl_rom_n_917, gl_rom_n_918, gl_rom_n_919, gl_rom_n_920, gl_rom_n_921 : std_logic;
  signal gl_rom_n_922, gl_rom_n_923, gl_rom_n_924, gl_rom_n_925, gl_rom_n_926 : std_logic;
  signal gl_rom_n_927, gl_rom_n_928, gl_rom_n_929, gl_rom_n_930, gl_rom_n_931 : std_logic;
  signal gl_rom_n_932, gl_rom_n_933, gl_rom_n_934, gl_rom_n_935, gl_rom_n_936 : std_logic;
  signal gl_rom_n_937, gl_rom_n_938, gl_rom_n_939, gl_rom_n_940, gl_rom_n_941 : std_logic;
  signal gl_rom_n_942, gl_rom_n_943, gl_rom_n_944, gl_rom_n_945, gl_rom_n_946 : std_logic;
  signal gl_rom_n_947, gl_rom_n_948, gl_rom_n_949, gl_rom_n_950, gl_rom_n_951 : std_logic;
  signal gl_rom_n_952, gl_rom_n_953, gl_rom_n_954, gl_rom_n_955, gl_rom_n_956 : std_logic;
  signal gl_rom_n_957, gl_rom_n_958, gl_rom_n_959, gl_rom_n_960, gl_rom_n_961 : std_logic;
  signal gl_rom_n_962, gl_rom_n_963, gl_rom_n_964, gl_rom_n_965, gl_rom_n_966 : std_logic;
  signal gl_rom_n_967, gl_rom_n_968, gl_rom_n_969, gl_rom_n_970, gl_rom_n_971 : std_logic;
  signal gl_rom_n_972, gl_rom_n_973, gl_rom_n_974, gl_rom_n_975, gl_rom_n_976 : std_logic;
  signal gl_rom_n_977, gl_rom_n_978, gl_rom_n_979, gl_rom_n_980, gl_rom_n_981 : std_logic;
  signal gl_rom_n_982, gl_rom_n_983, gl_rom_n_984, gl_rom_n_985, gl_rom_n_986 : std_logic;
  signal gl_rom_n_987, gl_rom_n_988, gl_rom_n_989, gl_rom_n_990, gl_rom_n_991 : std_logic;
  signal gl_rom_n_992, gl_rom_n_993, gl_rom_n_994, gl_rom_n_995, gl_rom_n_996 : std_logic;
  signal gl_rom_n_997, gl_rom_n_998, gl_rom_n_999, gl_rom_n_1000, gl_rom_n_1001 : std_logic;
  signal gl_rom_n_1002, gl_rom_n_1003, gl_rom_n_1004, gl_rom_n_1005, gl_rom_n_1006 : std_logic;
  signal gl_rom_n_1007, gl_rom_n_1008, gl_rom_n_1009, gl_rom_n_1010, gl_rom_n_1011 : std_logic;
  signal gl_rom_n_1012, gl_rom_n_1013, gl_rom_n_1014, gl_rom_n_1015, gl_rom_n_1016 : std_logic;
  signal gl_rom_n_1017, gl_rom_n_1018, gl_rom_n_1019, gl_rom_n_1020, gl_rom_n_1021 : std_logic;
  signal gl_rom_n_1022, gl_rom_n_1023, gl_rom_n_1024, gl_rom_n_1025, gl_rom_n_1026 : std_logic;
  signal gl_rom_n_1027, gl_rom_n_1028, gl_rom_n_1029, gl_rom_n_1030, gl_rom_n_1031 : std_logic;
  signal gl_rom_n_1032, gl_rom_n_1033, gl_rom_n_1034, gl_rom_n_1035, gl_rom_n_1036 : std_logic;
  signal gl_rom_n_1037, gl_rom_n_1038, gl_rom_n_1039, gl_rom_n_1040, gl_rom_n_1041 : std_logic;
  signal gl_rom_n_1042, gl_rom_n_1043, gl_rom_n_1044, gl_rom_n_1045, gl_rom_n_1046 : std_logic;
  signal gl_rom_n_1047, gl_rom_n_1048, gl_rom_n_1049, gl_rom_n_1050, gl_rom_n_1051 : std_logic;
  signal gl_rom_n_1052, gl_rom_n_1053, gl_rom_n_1054, gl_rom_n_1055, gl_rom_n_1056 : std_logic;
  signal gl_rom_n_1057, gl_rom_n_1058, gl_rom_n_1059, gl_rom_n_1060, gl_rom_n_1061 : std_logic;
  signal gl_rom_n_1062, gl_rom_n_1063, gl_rom_n_1064, gl_rom_n_1065, gl_rom_n_1066 : std_logic;
  signal gl_rom_n_1067, gl_rom_n_1068, gl_rom_n_1069, gl_rom_n_1070, gl_rom_n_1071 : std_logic;
  signal gl_rom_n_1072, gl_rom_n_1073, gl_rom_n_1074, gl_rom_n_1075, gl_rom_n_1076 : std_logic;
  signal gl_rom_n_1077, gl_rom_n_1078, gl_rom_n_1079, gl_rom_n_1080, gl_rom_n_1081 : std_logic;
  signal gl_rom_n_1082, gl_rom_n_1083, gl_rom_n_1084, gl_rom_n_1085, gl_rom_n_1086 : std_logic;
  signal gl_rom_n_1087, gl_rom_n_1088, gl_rom_n_1089, gl_rom_n_1090, gl_rom_n_1091 : std_logic;
  signal gl_rom_n_1092, gl_rom_n_1093, gl_rom_n_1094, gl_rom_n_1095, gl_rom_n_1096 : std_logic;
  signal gl_rom_n_1097, gl_rom_n_1098, gl_rom_n_1099, gl_rom_n_1100, gl_rom_n_1101 : std_logic;
  signal gl_rom_n_1102, gl_rom_n_1103, gl_rom_n_1104, gl_rom_n_1105, gl_rom_n_1106 : std_logic;
  signal gl_rom_n_1107, gl_rom_n_1108, gl_rom_n_1109, gl_rom_n_1110, gl_rom_n_1111 : std_logic;
  signal gl_rom_n_1112, gl_rom_n_1113, gl_rom_n_1114, gl_rom_n_1115, gl_rom_n_1116 : std_logic;
  signal gl_rom_n_1117, gl_rom_n_1118, gl_rom_n_1119, gl_rom_n_1120, gl_rom_n_1121 : std_logic;
  signal gl_rom_n_1122, gl_rom_n_1123, gl_rom_n_1124, gl_rom_n_1125, gl_rom_n_1126 : std_logic;
  signal gl_rom_n_1127, gl_rom_n_1128, gl_rom_n_1129, gl_rom_n_1130, gl_rom_n_1131 : std_logic;
  signal gl_rom_n_1132, gl_rom_n_1133, gl_rom_n_1134, gl_rom_n_1135, gl_rom_n_1136 : std_logic;
  signal gl_rom_n_1137, gl_rom_n_1138, gl_rom_n_1139, gl_rom_n_1140, gl_rom_n_1141 : std_logic;
  signal gl_rom_n_1142, gl_rom_n_1143, gl_rom_n_1144, gl_rom_n_1145, gl_rom_n_1146 : std_logic;
  signal gl_rom_n_1147, gl_rom_n_1148, gl_rom_n_1149, gl_rom_n_1150, gl_rom_n_1151 : std_logic;
  signal gl_rom_n_1152, gl_rom_n_1153, gl_rom_n_1154, gl_rom_n_1155, gl_rom_n_1156 : std_logic;
  signal gl_rom_n_1157, gl_rom_n_1158, gl_rom_n_1159, gl_rom_n_1160, gl_rom_n_1161 : std_logic;
  signal gl_rom_n_1162, gl_rom_n_1163, gl_rom_n_1164, gl_rom_n_1165, gl_rom_n_1166 : std_logic;
  signal gl_rom_n_1167, gl_rom_n_1168, gl_rom_n_1169, gl_rom_n_1170, gl_rom_n_1171 : std_logic;
  signal gl_rom_n_1172, gl_rom_n_1173, gl_rom_n_1174, gl_rom_n_1175, gl_rom_n_1176 : std_logic;
  signal gl_rom_n_1177, gl_rom_n_1178, gl_rom_n_1179, gl_rom_n_1180, gl_rom_n_1181 : std_logic;
  signal gl_rom_n_1182, gl_rom_n_1183, gl_rom_n_1184, gl_rom_n_1185, gl_rom_n_1186 : std_logic;
  signal gl_rom_n_1187, gl_rom_n_1188, gl_rom_n_1189, gl_rom_n_1190, gl_rom_n_1191 : std_logic;
  signal gl_rom_n_1192, gl_rom_n_1193, gl_rom_n_1194, gl_rom_n_1195, gl_rom_n_1196 : std_logic;
  signal gl_rom_n_1197, gl_rom_n_1198, gl_rom_n_1199, gl_rom_n_1200, gl_rom_n_1201 : std_logic;
  signal gl_rom_n_1202, gl_rom_n_1203, gl_rom_n_1204, gl_rom_n_1205, gl_rom_n_1206 : std_logic;
  signal gl_rom_n_1207, gl_rom_n_1208, gl_rom_n_1209, gl_rom_n_1210, gl_rom_n_1211 : std_logic;
  signal gl_rom_n_1212, gl_rom_n_1213, gl_rom_n_1214, gl_rom_n_1215, gl_rom_n_1216 : std_logic;
  signal gl_rom_n_1217, gl_rom_n_1218, gl_rom_n_1219, gl_rom_n_1220, gl_rom_n_1221 : std_logic;
  signal gl_rom_n_1222, gl_rom_n_1223, gl_rom_n_1224, gl_rom_n_1225, gl_rom_n_1226 : std_logic;
  signal gl_rom_n_1227, gl_rom_n_1228, gl_rom_n_1229, gl_rom_n_1230, gl_rom_n_1231 : std_logic;
  signal gl_rom_n_1232, gl_rom_n_1233, gl_rom_n_1234, gl_rom_n_1235, gl_rom_n_1236 : std_logic;
  signal gl_rom_n_1237, gl_rom_n_1238, gl_rom_n_1239, gl_rom_n_1240, gl_rom_n_1241 : std_logic;
  signal gl_rom_n_1242, gl_rom_n_1243, gl_rom_n_1244, gl_rom_n_1245, gl_rom_n_1246 : std_logic;
  signal gl_rom_n_1247, gl_rom_n_1248, gl_rom_n_1249, gl_rom_n_1250, gl_rom_n_1251 : std_logic;
  signal gl_rom_n_1252, gl_rom_n_1253, gl_rom_n_1254, gl_rom_n_1255, gl_rom_n_1256 : std_logic;
  signal gl_rom_n_1257, gl_rom_n_1258, gl_rom_n_1259, gl_rom_n_1260, gl_rom_n_1261 : std_logic;
  signal gl_rom_n_1262, gl_rom_n_1263, gl_rom_n_1264, gl_rom_n_1265, gl_rom_n_1266 : std_logic;
  signal gl_rom_n_1267, gl_rom_n_1268, gl_rom_n_1269, gl_rom_n_1270, gl_rom_n_1271 : std_logic;
  signal gl_rom_n_1272, gl_rom_n_1273, gl_rom_n_1274, gl_rom_n_1275, gl_rom_n_1276 : std_logic;
  signal gl_rom_n_1277, gl_rom_n_1278, gl_rom_n_1279, gl_rom_n_1280, gl_rom_n_1281 : std_logic;
  signal gl_rom_n_1282, gl_rom_n_1283, gl_rom_n_1284, gl_rom_n_1285, gl_rom_n_1286 : std_logic;
  signal gl_rom_n_1287, gl_rom_n_1288, gl_rom_n_1289, gl_rom_n_1290, gl_rom_n_1291 : std_logic;
  signal gl_rom_n_1292, gl_rom_n_1293, gl_rom_n_1294, gl_rom_n_1295, gl_rom_n_1296 : std_logic;
  signal gl_rom_n_1297, gl_rom_n_1298, gl_rom_n_1299, gl_rom_n_1300, gl_rom_n_1301 : std_logic;
  signal gl_rom_n_1302, gl_rom_n_1303, gl_rom_n_1304, gl_rom_n_1305, gl_rom_n_1306 : std_logic;
  signal gl_rom_n_1307, gl_rom_n_1308, gl_rom_n_1309, gl_rom_n_1310, gl_rom_n_1311 : std_logic;
  signal gl_rom_n_1312, gl_rom_n_1313, gl_rom_n_1314, gl_rom_n_1315, gl_rom_n_1316 : std_logic;
  signal gl_rom_n_1317, gl_rom_n_1318, gl_rom_n_1319, gl_rom_n_1320, gl_rom_n_1321 : std_logic;
  signal gl_rom_n_1322, gl_rom_n_1323, gl_rom_n_1324, gl_rom_n_1325, gl_rom_n_1326 : std_logic;
  signal gl_rom_n_1327, gl_rom_n_1328, gl_rom_n_1329, gl_rom_n_1330, gl_rom_n_1331 : std_logic;
  signal gl_rom_n_1332, gl_rom_n_1333, gl_rom_n_1334, gl_rom_n_1335, gl_rom_n_1336 : std_logic;
  signal gl_rom_n_1337, gl_rom_n_1338, gl_rom_n_1339, gl_rom_n_1340, gl_rom_n_1341 : std_logic;
  signal gl_rom_n_1342, gl_rom_n_1343, gl_rom_n_1344, gl_rom_n_1345, gl_rom_n_1346 : std_logic;
  signal gl_rom_n_1347, gl_rom_n_1348, gl_rom_n_1349, gl_rom_n_1350, gl_rom_n_1351 : std_logic;
  signal gl_rom_n_1352, gl_rom_n_1353, gl_rom_n_1354, gl_rom_n_1355, gl_rom_n_1356 : std_logic;
  signal gl_rom_n_1357, gl_rom_n_1358, gl_rom_n_1359, gl_rom_n_1360, gl_rom_n_1361 : std_logic;
  signal gl_rom_n_1362, gl_rom_n_1363, gl_rom_n_1364, gl_rom_n_1365, gl_rom_n_1366 : std_logic;
  signal gl_rom_n_1367, gl_rom_n_1368, gl_rom_n_1369, gl_rom_n_1370, gl_rom_n_1371 : std_logic;
  signal gl_rom_n_1372, gl_rom_n_1373, gl_rom_n_1374, gl_rom_n_1375, gl_rom_n_1376 : std_logic;
  signal gl_rom_n_1377, gl_rom_n_1378, gl_rom_n_1379, gl_rom_n_1380, gl_rom_n_1381 : std_logic;
  signal gl_rom_n_1382, gl_rom_n_1383, gl_rom_n_1384, gl_rom_n_1385, gl_rom_n_1386 : std_logic;
  signal gl_rom_n_1387, gl_rom_n_1388, gl_rom_n_1389, gl_rom_n_1390, gl_rom_n_1391 : std_logic;
  signal gl_rom_n_1392, gl_rom_n_1393, gl_rom_n_1394, gl_rom_n_1395, gl_rom_n_1396 : std_logic;
  signal gl_rom_n_1397, gl_rom_n_1398, gl_rom_n_1399, gl_rom_n_1400, gl_rom_n_1401 : std_logic;
  signal gl_rom_n_1402, gl_rom_n_1403, gl_rom_n_1404, gl_rom_n_1405, gl_rom_n_1406 : std_logic;
  signal gl_rom_n_1407, gl_rom_n_1408, gl_rom_n_1409, gl_rom_n_1410, gl_rom_n_1411 : std_logic;
  signal gl_rom_n_1412, gl_rom_n_1413, gl_rom_n_1414, gl_rom_n_1415, gl_rom_n_1416 : std_logic;
  signal gl_rom_n_1417, gl_rom_n_1418, gl_rom_n_1419, gl_rom_n_1420, gl_rom_n_1421 : std_logic;
  signal gl_rom_n_1422, gl_rom_n_1423, gl_rom_n_1424, gl_rom_n_1425, gl_rom_n_1426 : std_logic;
  signal gl_rom_n_1427, gl_rom_n_1428, gl_rom_n_1429, gl_rom_n_1430, gl_rom_n_1431 : std_logic;
  signal gl_rom_n_1432, gl_rom_n_1433, gl_rom_n_1434, gl_rom_n_1435, gl_rom_n_1436 : std_logic;
  signal gl_rom_n_1437, gl_rom_n_1438, gl_rom_n_1439, gl_rom_n_1440, gl_rom_n_1441 : std_logic;
  signal gl_rom_n_1442, gl_rom_n_1443, gl_rom_n_1444, gl_rom_n_1445, gl_rom_n_1446 : std_logic;
  signal gl_rom_n_1447, gl_rom_n_1448, gl_rom_n_1449, gl_rom_n_1450, gl_rom_n_1451 : std_logic;
  signal gl_rom_n_1452, gl_rom_n_1453, gl_rom_n_1454, gl_rom_n_1455, gl_rom_n_1456 : std_logic;
  signal gl_rom_n_1457, gl_rom_n_1458, gl_rom_n_1459, gl_rom_n_1460, gl_rom_n_1461 : std_logic;
  signal gl_rom_n_1462, gl_rom_n_1463, gl_rom_n_1464, gl_rom_n_1465, gl_rom_n_1466 : std_logic;
  signal gl_rom_n_1467, gl_rom_n_1468, gl_rom_n_1469, gl_rom_n_1470, gl_rom_n_1471 : std_logic;
  signal gl_rom_n_1472, gl_rom_n_1473, gl_rom_n_1474, gl_rom_n_1475, gl_rom_n_1476 : std_logic;
  signal gl_rom_n_1477, gl_rom_n_1478, gl_rom_n_1479, gl_rom_n_1480, gl_rom_n_1481 : std_logic;
  signal gl_rom_n_1482, gl_rom_n_1483, gl_rom_n_1484, gl_rom_n_1485, gl_rom_n_1486 : std_logic;
  signal gl_rom_n_1487, gl_rom_n_1488, gl_rom_n_1489, gl_rom_n_1490, gl_rom_n_1491 : std_logic;
  signal gl_rom_n_1492, gl_rom_n_1493, gl_rom_n_1494, gl_rom_n_1495, gl_rom_n_1496 : std_logic;
  signal gl_rom_n_1497, gl_rom_n_1498, gl_rom_n_1499, gl_rom_n_1500, gl_sig_blue : std_logic;
  signal gl_sig_countdown_aan, gl_sig_green, gl_sig_red, gl_sig_scale_h, gl_sig_scale_v : std_logic;
  signal gl_vgd_n_0, gl_vgd_n_1, gl_vgd_n_2, gl_vgd_n_3, gl_vgd_n_4 : std_logic;
  signal gl_vgd_n_5, gl_vgd_n_6, gl_vgd_n_7, gl_vgd_n_8, gl_vgd_n_9 : std_logic;
  signal gl_vgd_n_10, gl_vgd_n_11, gl_vgd_n_12, gl_vgd_n_13, gl_vgd_n_14 : std_logic;
  signal gl_vgd_n_15, gl_vgd_n_16, gl_vgd_n_17, gl_vgd_n_18, gl_vgd_n_19 : std_logic;
  signal gl_vgd_n_20, gl_vgd_n_21, gl_vgd_n_22, gl_vgd_n_23, gl_vgd_n_24 : std_logic;
  signal gl_vgd_n_25, gl_vgd_n_26, gl_vgd_n_27, gl_vgd_n_28, gl_vgd_n_29 : std_logic;
  signal gl_vgd_n_30, gl_vgd_n_31, gl_vgd_n_32, gl_vgd_n_33, gl_vgd_n_34 : std_logic;
  signal gl_vgd_n_35, gl_vgd_n_36, gl_vgd_n_37, gl_vgd_n_38, gl_vgd_n_39 : std_logic;
  signal gl_vgd_n_40, gl_vgd_n_41, gl_vgd_n_42, gl_vgd_n_43, gl_vgd_n_44 : std_logic;
  signal gl_vgd_n_45, gl_vgd_n_46, gl_vgd_n_47, gl_vgd_n_48, gl_vgd_n_49 : std_logic;
  signal gl_vgd_n_50, gl_vgd_n_51, gl_vgd_n_52, gl_vgd_n_53, gl_vgd_n_54 : std_logic;
  signal gl_vgd_n_55, gl_vgd_n_56, gl_vgd_n_57, gl_vgd_n_58, gl_vgd_n_59 : std_logic;
  signal gl_vgd_n_60, gl_vgd_n_61, gl_vgd_n_62, gl_vgd_n_63, gl_vgd_n_64 : std_logic;
  signal gl_vgd_n_65, gl_vgd_n_67, gl_vgd_n_68, gl_vgd_n_69, gl_vgd_n_70 : std_logic;
  signal gl_vgd_n_71, gl_vgd_n_72, gl_vgd_n_73, gl_vgd_n_74, gl_vgd_n_75 : std_logic;
  signal gl_vgd_n_76, gl_vgd_n_77, gl_vgd_n_78, gl_vgd_n_79, gl_vgd_n_80 : std_logic;
  signal gl_vgd_n_81, ml_handshake_mouse_out, ml_il_color1_n_0, ml_il_color1_n_1, ml_il_color1_n_2 : std_logic;
  signal ml_il_color1_n_3, ml_il_color1_n_4, ml_il_color1_n_5, ml_il_color1_n_6, ml_il_color1_n_7 : std_logic;
  signal ml_il_color1_n_8, ml_il_color1_n_9, ml_il_color1_n_10, ml_il_color1_n_11, ml_il_color1_n_12 : std_logic;
  signal ml_il_color1_n_13, ml_il_color1_n_14, ml_il_color1_n_15, ml_il_color1_n_16, ml_il_color1_n_17 : std_logic;
  signal ml_il_color1_n_22, ml_il_color1_n_23, ml_il_x1_n_0, ml_il_x1_n_1, ml_il_x1_n_2 : std_logic;
  signal ml_il_x1_n_3, ml_il_x1_n_4, ml_il_x1_n_5, ml_il_x1_n_6, ml_il_x1_n_7 : std_logic;
  signal ml_il_x1_n_8, ml_il_x1_n_9, ml_il_x1_n_10, ml_il_x1_n_11, ml_il_x1_n_12 : std_logic;
  signal ml_il_x1_n_13, ml_il_x1_n_14, ml_il_x1_n_15, ml_il_x1_n_16, ml_il_x1_n_17 : std_logic;
  signal ml_il_x1_n_18, ml_il_x1_n_19, ml_il_x1_n_20, ml_il_x1_n_21, ml_il_x1_n_22 : std_logic;
  signal ml_il_x1_n_23, ml_il_x1_n_24, ml_il_x1_n_25, ml_il_x1_n_26, ml_il_x1_n_27 : std_logic;
  signal ml_il_x1_n_28, ml_il_x1_n_29, ml_il_y1_n_0, ml_il_y1_n_1, ml_il_y1_n_2 : std_logic;
  signal ml_il_y1_n_3, ml_il_y1_n_4, ml_il_y1_n_5, ml_il_y1_n_7, ml_il_y1_n_8 : std_logic;
  signal ml_il_y1_n_9, ml_il_y1_n_10, ml_il_y1_n_11, ml_il_y1_n_12, ml_il_y1_n_13 : std_logic;
  signal ml_il_y1_n_14, ml_il_y1_n_17, ml_il_y1_n_18, ml_il_y1_n_20, ml_il_y1_n_22 : std_logic;
  signal ml_il_y1_n_23, ml_il_y1_n_24, ml_il_y1_n_25, ml_il_y1_n_26, ml_il_y1_n_27 : std_logic;
  signal ml_il_y1_n_28, ml_il_y1_n_29, ml_il_y1_n_30, ml_il_y1_n_31, ml_il_y1_n_32 : std_logic;
  signal ml_il_y1_n_33, ml_il_y1_n_36, ml_il_y1_n_39, ml_il_y1_n_40, ml_il_y1_n_41 : std_logic;
  signal ml_ms_Clk15k_buffered, ml_ms_Clk15k_intermediate, ml_ms_Data_in_buffered, ml_ms_Data_in_intermediate, ml_ms_actBit : std_logic;
  signal ml_ms_btnflipfloprst, ml_ms_cntD_n_0, ml_ms_cntD_n_1, ml_ms_cntD_n_2, ml_ms_cntD_n_3 : std_logic;
  signal ml_ms_cntD_n_4, ml_ms_cntD_n_5, ml_ms_cntD_n_6, ml_ms_cntD_n_7, ml_ms_cntD_n_8 : std_logic;
  signal ml_ms_cntD_n_9, ml_ms_cntD_n_10, ml_ms_cntD_n_11, ml_ms_cntD_n_12, ml_ms_cntD_n_13 : std_logic;
  signal ml_ms_cntD_n_14, ml_ms_cntD_n_15, ml_ms_cntD_n_16, ml_ms_cntD_n_17, ml_ms_cntD_n_18 : std_logic;
  signal ml_ms_cntD_n_19, ml_ms_cntD_n_20, ml_ms_cntD_n_21, ml_ms_cntD_n_22, ml_ms_cntD_n_23 : std_logic;
  signal ml_ms_cntReset15K, ml_ms_cntReset25M, ml_ms_cntReset25M_main, ml_ms_cntReset25M_send, ml_ms_cnt_n_0 : std_logic;
  signal ml_ms_cnt_n_1, ml_ms_cnt_n_2, ml_ms_cnt_n_3, ml_ms_cnt_n_4, ml_ms_cnt_n_5 : std_logic;
  signal ml_ms_cnt_n_6, ml_ms_cnt_n_7, ml_ms_cnt_n_8, ml_ms_cnt_n_9, ml_ms_cnt_n_10 : std_logic;
  signal ml_ms_cnt_n_11, ml_ms_cnt_n_12, ml_ms_cnt_n_13, ml_ms_cnt_n_14, ml_ms_cnt_n_15 : std_logic;
  signal ml_ms_cnt_n_16, ml_ms_cnt_n_17, ml_ms_cnt_n_18, ml_ms_cnt_n_19, ml_ms_cnt_n_20 : std_logic;
  signal ml_ms_cnt_n_21, ml_ms_cnt_n_22, ml_ms_cnt_n_23, ml_ms_count_debounce_reset, ml_ms_ed_n_0 : std_logic;
  signal ml_ms_ed_n_1, ml_ms_ed_n_2, ml_ms_ed_n_3, ml_ms_ed_n_4, ml_ms_ed_n_5 : std_logic;
  signal ml_ms_ed_n_6, ml_ms_ed_n_7, ml_ms_ed_n_8, ml_ms_ed_n_9, ml_ms_ed_n_10 : std_logic;
  signal ml_ms_ed_n_12, ml_ms_ed_n_13, ml_ms_ed_n_14, ml_ms_ed_n_15, ml_ms_ed_n_16 : std_logic;
  signal ml_ms_ed_n_35, ml_ms_ed_reg1, ml_ms_ed_reg2, ml_ms_flipflop1_Q_9, ml_ms_flipflop4_Q_9 : std_logic;
  signal ml_ms_flipflop5_Q_9, ml_ms_flipflop6_Q_9, ml_ms_mfsm_n_0, ml_ms_mfsm_n_1, ml_ms_mfsm_n_2 : std_logic;
  signal ml_ms_mfsm_n_3, ml_ms_mfsm_n_4, ml_ms_mfsm_n_5, ml_ms_mfsm_n_6, ml_ms_mfsm_n_7 : std_logic;
  signal ml_ms_mfsm_n_8, ml_ms_mfsm_n_9, ml_ms_mfsm_n_10, ml_ms_mfsm_n_11, ml_ms_mfsm_n_12 : std_logic;
  signal ml_ms_mfsm_n_13, ml_ms_mfsm_n_14, ml_ms_mfsm_n_15, ml_ms_mfsm_n_16, ml_ms_mfsm_n_17 : std_logic;
  signal ml_ms_mfsm_n_18, ml_ms_mfsm_n_19, ml_ms_mfsm_n_20, ml_ms_mfsm_n_21, ml_ms_mfsm_n_22 : std_logic;
  signal ml_ms_mfsm_n_23, ml_ms_mfsm_n_24, ml_ms_mfsm_n_25, ml_ms_mfsm_n_26, ml_ms_mfsm_n_27 : std_logic;
  signal ml_ms_mfsm_n_28, ml_ms_mfsm_n_29, ml_ms_mfsm_n_30, ml_ms_mfsm_n_31, ml_ms_mfsm_n_32 : std_logic;
  signal ml_ms_mfsm_n_33, ml_ms_mfsm_n_34, ml_ms_mfsm_n_35, ml_ms_mfsm_n_36, ml_ms_mfsm_n_37 : std_logic;
  signal ml_ms_mfsm_n_38, ml_ms_mfsm_n_39, ml_ms_mfsm_n_40, ml_ms_mfsm_n_41, ml_ms_mfsm_n_43 : std_logic;
  signal ml_ms_mfsm_n_45, ml_ms_mfsm_n_46, ml_ms_mfsm_n_47, ml_ms_mfsm_n_48, ml_ms_mfsm_n_49 : std_logic;
  signal ml_ms_mfsm_n_50, ml_ms_mfsm_n_51, ml_ms_mfsm_n_52, ml_ms_mfsm_n_53, ml_ms_mfsm_n_54 : std_logic;
  signal ml_ms_mfsm_n_55, ml_ms_mfsm_n_56, ml_ms_mfsm_n_57, ml_ms_mfsm_n_58, ml_ms_mfsm_n_59 : std_logic;
  signal ml_ms_mfsm_n_60, ml_ms_mfsm_n_61, ml_ms_mfsm_n_62, ml_ms_mfsm_n_63, ml_ms_mfsm_n_64 : std_logic;
  signal ml_ms_mfsm_n_65, ml_ms_mfsm_n_66, ml_ms_mfsm_n_67, ml_ms_mfsm_n_68, ml_ms_mfsm_n_69 : std_logic;
  signal ml_ms_mfsm_n_70, ml_ms_mfsm_n_71, ml_ms_mfsm_n_72, ml_ms_mfsm_n_73, ml_ms_mfsm_n_74 : std_logic;
  signal ml_ms_mfsm_n_75, ml_ms_mfsm_n_148, ml_ms_muxFSM, ml_ms_muxReg, ml_ms_mux_select : std_logic;
  signal ml_ms_mux_select_main, ml_ms_mx_n_0, ml_ms_mx_n_1, ml_ms_n_0, ml_ms_n_1 : std_logic;
  signal ml_ms_n_2, ml_ms_n_3, ml_ms_n_4, ml_ms_n_5, ml_ms_n_6 : std_logic;
  signal ml_ms_n_7, ml_ms_n_8, ml_ms_n_9, ml_ms_n_10, ml_ms_n_11 : std_logic;
  signal ml_ms_n_12, ml_ms_n_13, ml_ms_n_14, ml_ms_n_15, ml_ms_n_16 : std_logic;
  signal ml_ms_n_17, ml_ms_n_18, ml_ms_n_19, ml_ms_n_20, ml_ms_n_21 : std_logic;
  signal ml_ms_n_22, ml_ms_n_23, ml_ms_n_24, ml_ms_n_25, ml_ms_n_26 : std_logic;
  signal ml_ms_n_27, ml_ms_n_28, ml_ms_n_29, ml_ms_n_30, ml_ms_n_31 : std_logic;
  signal ml_ms_n_32, ml_ms_n_33, ml_ms_n_34, ml_ms_n_35, ml_ms_n_36 : std_logic;
  signal ml_ms_n_37, ml_ms_n_38, ml_ms_n_39, ml_ms_n_40, ml_ms_n_41 : std_logic;
  signal ml_ms_n_42, ml_ms_n_43, ml_ms_n_44, ml_ms_n_45, ml_ms_n_46 : std_logic;
  signal ml_ms_n_47, ml_ms_n_48, ml_ms_n_49, ml_ms_n_50, ml_ms_n_51 : std_logic;
  signal ml_ms_n_52, ml_ms_n_53, ml_ms_n_54, ml_ms_n_55, ml_ms_n_56 : std_logic;
  signal ml_ms_n_57, ml_ms_n_58, ml_ms_n_59, ml_ms_n_60, ml_ms_n_61 : std_logic;
  signal ml_ms_n_62, ml_ms_n_63, ml_ms_n_78, ml_ms_n_82, ml_ms_output_edgedet : std_logic;
  signal ml_ms_reset_send, ml_ms_sfsm_n_383, ml_ms_sr11_data_out_0_79, ml_ms_sr11_data_out_1_80, ml_ms_sr11_data_out_2_81 : std_logic;
  signal ml_ms_sr11_data_out_3_82, ml_ms_sr11_n_0, ml_ms_tb_n_0, ml_ms_tb_n_1, ml_ms_tb_n_2 : std_logic;
  signal ml_ms_tb_n_3, ml_ms_tb_n_4, ml_ms_tb_n_5, ml_ms_tb_n_6, ml_ms_timerReset : std_logic;
  signal ml_ms_xflipfloprst, ml_ms_yflipfloprst, n_0, sig_draw, sig_middelsteknop : std_logic;

begin

  ml_ms_timr : mouse_timer port map(clk => clk, reset => ml_ms_timerReset, count_out => ml_ms_timer_count);
  g1 : BUFFD4BWP7T port map(I => reset, Z => n_0);
  gl_rom_rom_colour_out_reg_0 : LHQD1BWP7T port map(E => clk, D => gl_rom_n_1500, Q => gl_sig_rom(0));
  gl_rom_rom_colour_out_reg_1 : LHQD1BWP7T port map(E => clk, D => gl_rom_n_1499, Q => gl_sig_rom(1));
  gl_rom_g34920 : MOAI22D0BWP7T port map(A1 => gl_rom_n_1496, A2 => gl_sig_e(9), B1 => gl_rom_n_1498, B2 => gl_sig_e(9), ZN => gl_rom_n_1500);
  gl_rom_g34921 : MOAI22D0BWP7T port map(A1 => gl_rom_n_1497, A2 => gl_sig_e(9), B1 => gl_rom_n_1495, B2 => gl_sig_e(9), ZN => gl_rom_n_1499);
  gl_rom_g34922 : ND4D0BWP7T port map(A1 => gl_rom_n_1481, A2 => gl_rom_n_1490, A3 => gl_rom_n_1480, A4 => gl_rom_n_1488, ZN => gl_rom_n_1498);
  gl_rom_g34923 : AN4D0BWP7T port map(A1 => gl_rom_n_1482, A2 => gl_rom_n_1483, A3 => gl_rom_n_1484, A4 => gl_rom_n_1493, Z => gl_rom_n_1497);
  gl_rom_g34924 : AN4D0BWP7T port map(A1 => gl_rom_n_1494, A2 => gl_rom_n_1485, A3 => gl_rom_n_1487, A4 => gl_rom_n_1492, Z => gl_rom_n_1496);
  gl_rom_g34925 : ND4D0BWP7T port map(A1 => gl_rom_n_1489, A2 => gl_rom_n_1491, A3 => gl_rom_n_1486, A4 => gl_rom_n_1479, ZN => gl_rom_n_1495);
  gl_rom_g34926 : AOI22D0BWP7T port map(A1 => gl_rom_n_1475, A2 => gl_rom_n_33, B1 => gl_rom_n_1463, B2 => gl_rom_n_36, ZN => gl_rom_n_1494);
  gl_rom_g34927 : AOI22D0BWP7T port map(A1 => gl_rom_n_1472, A2 => gl_rom_n_37, B1 => gl_rom_n_1456, B2 => gl_rom_n_31, ZN => gl_rom_n_1493);
  gl_rom_g34928 : AOI22D0BWP7T port map(A1 => gl_rom_n_1460, A2 => gl_rom_n_37, B1 => gl_rom_n_1447, B2 => gl_rom_n_31, ZN => gl_rom_n_1492);
  gl_rom_g34929 : AOI22D0BWP7T port map(A1 => gl_rom_n_1477, A2 => gl_rom_n_37, B1 => gl_rom_n_1462, B2 => gl_rom_n_31, ZN => gl_rom_n_1491);
  gl_rom_g34930 : AOI22D0BWP7T port map(A1 => gl_rom_n_1458, A2 => gl_rom_n_37, B1 => gl_rom_n_1454, B2 => gl_rom_n_31, ZN => gl_rom_n_1490);
  gl_rom_g34931 : AOI22D0BWP7T port map(A1 => gl_rom_n_1474, A2 => gl_rom_n_32, B1 => gl_rom_n_1476, B2 => gl_rom_n_35, ZN => gl_rom_n_1489);
  gl_rom_g34932 : AOI22D0BWP7T port map(A1 => gl_rom_n_1452, A2 => gl_rom_n_32, B1 => gl_rom_n_1473, B2 => gl_rom_n_35, ZN => gl_rom_n_1488);
  gl_rom_g34933 : AOI22D0BWP7T port map(A1 => gl_rom_n_1470, A2 => gl_rom_n_38, B1 => gl_rom_n_1455, B2 => gl_rom_n_34, ZN => gl_rom_n_1487);
  gl_rom_g34934 : AOI22D0BWP7T port map(A1 => gl_rom_n_1449, A2 => gl_rom_n_33, B1 => gl_rom_n_1478, B2 => gl_rom_n_36, ZN => gl_rom_n_1486);
  gl_rom_g34935 : AOI22D0BWP7T port map(A1 => gl_rom_n_1465, A2 => gl_rom_n_32, B1 => gl_rom_n_1467, B2 => gl_rom_n_35, ZN => gl_rom_n_1485);
  gl_rom_g34936 : AOI22D0BWP7T port map(A1 => gl_rom_n_1466, A2 => gl_rom_n_33, B1 => gl_rom_n_1453, B2 => gl_rom_n_36, ZN => gl_rom_n_1484);
  gl_rom_g34937 : AOI22D0BWP7T port map(A1 => gl_rom_n_1464, A2 => gl_rom_n_32, B1 => gl_rom_n_1451, B2 => gl_rom_n_35, ZN => gl_rom_n_1483);
  gl_rom_g34938 : AOI22D0BWP7T port map(A1 => gl_rom_n_1468, A2 => gl_rom_n_38, B1 => gl_rom_n_1469, B2 => gl_rom_n_34, ZN => gl_rom_n_1482);
  gl_rom_g34939 : AOI22D0BWP7T port map(A1 => gl_rom_n_1471, A2 => gl_rom_n_33, B1 => gl_rom_n_1448, B2 => gl_rom_n_36, ZN => gl_rom_n_1481);
  gl_rom_g34940 : AOI22D0BWP7T port map(A1 => gl_rom_n_1457, A2 => gl_rom_n_38, B1 => gl_rom_n_1450, B2 => gl_rom_n_34, ZN => gl_rom_n_1480);
  gl_rom_g34941 : AOI22D0BWP7T port map(A1 => gl_rom_n_1459, A2 => gl_rom_n_38, B1 => gl_rom_n_1461, B2 => gl_rom_n_34, ZN => gl_rom_n_1479);
  gl_rom_g34942 : ND4D0BWP7T port map(A1 => gl_rom_n_1342, A2 => gl_rom_n_1340, A3 => gl_rom_n_1424, A4 => gl_rom_n_1337, ZN => gl_rom_n_1478);
  gl_rom_g34943 : ND4D0BWP7T port map(A1 => gl_rom_n_1407, A2 => gl_rom_n_1409, A3 => gl_rom_n_1445, A4 => gl_rom_n_1404, ZN => gl_rom_n_1477);
  gl_rom_g34944 : ND4D0BWP7T port map(A1 => gl_rom_n_1403, A2 => gl_rom_n_1400, A3 => gl_rom_n_1398, A4 => gl_rom_n_1443, ZN => gl_rom_n_1476);
  gl_rom_g34945 : ND4D0BWP7T port map(A1 => gl_rom_n_1401, A2 => gl_rom_n_1392, A3 => gl_rom_n_1396, A4 => gl_rom_n_1442, ZN => gl_rom_n_1475);
  gl_rom_g34946 : ND4D0BWP7T port map(A1 => gl_rom_n_1397, A2 => gl_rom_n_1440, A3 => gl_rom_n_1391, A4 => gl_rom_n_1394, ZN => gl_rom_n_1474);
  gl_rom_g34947 : ND4D0BWP7T port map(A1 => gl_rom_n_1386, A2 => gl_rom_n_1366, A3 => gl_rom_n_1435, A4 => gl_rom_n_1381, ZN => gl_rom_n_1473);
  gl_rom_g34948 : ND4D0BWP7T port map(A1 => gl_rom_n_1385, A2 => gl_rom_n_1383, A3 => gl_rom_n_1379, A4 => gl_rom_n_1437, ZN => gl_rom_n_1472);
  gl_rom_g34949 : ND4D0BWP7T port map(A1 => gl_rom_n_1371, A2 => gl_rom_n_1427, A3 => gl_rom_n_1341, A4 => gl_rom_n_1350, ZN => gl_rom_n_1471);
  gl_rom_g34950 : ND4D0BWP7T port map(A1 => gl_rom_n_1377, A2 => gl_rom_n_1376, A3 => gl_rom_n_1434, A4 => gl_rom_n_1368, ZN => gl_rom_n_1470);
  gl_rom_g34951 : ND4D0BWP7T port map(A1 => gl_rom_n_1378, A2 => gl_rom_n_1436, A3 => gl_rom_n_1375, A4 => gl_rom_n_1374, ZN => gl_rom_n_1469);
  gl_rom_g34952 : ND4D0BWP7T port map(A1 => gl_rom_n_1372, A2 => gl_rom_n_1433, A3 => gl_rom_n_1369, A4 => gl_rom_n_1370, ZN => gl_rom_n_1468);
  gl_rom_g34953 : ND4D0BWP7T port map(A1 => gl_rom_n_1365, A2 => gl_rom_n_1357, A3 => gl_rom_n_1430, A4 => gl_rom_n_1363, ZN => gl_rom_n_1467);
  gl_rom_g34954 : ND4D0BWP7T port map(A1 => gl_rom_n_1359, A2 => gl_rom_n_1360, A3 => gl_rom_n_1429, A4 => gl_rom_n_1356, ZN => gl_rom_n_1466);
  gl_rom_g34955 : ND4D0BWP7T port map(A1 => gl_rom_n_1355, A2 => gl_rom_n_1347, A3 => gl_rom_n_1344, A4 => gl_rom_n_1426, ZN => gl_rom_n_1465);
  gl_rom_g34956 : ND4D0BWP7T port map(A1 => gl_rom_n_1348, A2 => gl_rom_n_1425, A3 => gl_rom_n_1346, A4 => gl_rom_n_1343, ZN => gl_rom_n_1464);
  gl_rom_g34957 : ND4D0BWP7T port map(A1 => gl_rom_n_1446, A2 => gl_rom_n_1405, A3 => gl_rom_n_1408, A4 => gl_rom_n_1414, ZN => gl_rom_n_1463);
  gl_rom_g34958 : ND4D0BWP7T port map(A1 => gl_rom_n_1415, A2 => gl_rom_n_1413, A3 => gl_rom_n_1412, A4 => gl_rom_n_1410, ZN => gl_rom_n_1462);
  gl_rom_g34959 : ND4D0BWP7T port map(A1 => gl_rom_n_1330, A2 => gl_rom_n_1325, A3 => gl_rom_n_1419, A4 => gl_rom_n_1327, ZN => gl_rom_n_1461);
  gl_rom_g34960 : ND4D0BWP7T port map(A1 => gl_rom_n_1329, A2 => gl_rom_n_1326, A3 => gl_rom_n_1418, A4 => gl_rom_n_1320, ZN => gl_rom_n_1460);
  gl_rom_g34961 : ND4D0BWP7T port map(A1 => gl_rom_n_1323, A2 => gl_rom_n_1417, A3 => gl_rom_n_1319, A4 => gl_rom_n_1324, ZN => gl_rom_n_1459);
  gl_rom_g34962 : ND4D0BWP7T port map(A1 => gl_rom_n_1441, A2 => gl_rom_n_1351, A3 => gl_rom_n_1373, A4 => gl_rom_n_1322, ZN => gl_rom_n_1458);
  gl_rom_g34963 : ND4D0BWP7T port map(A1 => gl_rom_n_1444, A2 => gl_rom_n_1399, A3 => gl_rom_n_1411, A4 => gl_rom_n_1393, ZN => gl_rom_n_1457);
  gl_rom_g34964 : ND4D0BWP7T port map(A1 => gl_rom_n_1388, A2 => gl_rom_n_1439, A3 => gl_rom_n_1390, A4 => gl_rom_n_1387, ZN => gl_rom_n_1456);
  gl_rom_g34965 : ND4D0BWP7T port map(A1 => gl_rom_n_1389, A2 => gl_rom_n_1438, A3 => gl_rom_n_1384, A4 => gl_rom_n_1380, ZN => gl_rom_n_1455);
  gl_rom_g34966 : ND4D0BWP7T port map(A1 => gl_rom_n_1402, A2 => gl_rom_n_1353, A3 => gl_rom_n_1361, A4 => gl_rom_n_1423, ZN => gl_rom_n_1454);
  gl_rom_g34967 : ND4D0BWP7T port map(A1 => gl_rom_n_1432, A2 => gl_rom_n_1362, A3 => gl_rom_n_1367, A4 => gl_rom_n_1364, ZN => gl_rom_n_1453);
  gl_rom_g34968 : ND4D0BWP7T port map(A1 => gl_rom_n_1431, A2 => gl_rom_n_1345, A3 => gl_rom_n_1358, A4 => gl_rom_n_1382, ZN => gl_rom_n_1452);
  gl_rom_g34969 : ND4D0BWP7T port map(A1 => gl_rom_n_1354, A2 => gl_rom_n_1428, A3 => gl_rom_n_1352, A4 => gl_rom_n_1349, ZN => gl_rom_n_1451);
  gl_rom_g34970 : ND4D0BWP7T port map(A1 => gl_rom_n_1333, A2 => gl_rom_n_1422, A3 => gl_rom_n_1328, A4 => gl_rom_n_1321, ZN => gl_rom_n_1450);
  gl_rom_g34971 : ND4D0BWP7T port map(A1 => gl_rom_n_1336, A2 => gl_rom_n_1335, A3 => gl_rom_n_1331, A4 => gl_rom_n_1421, ZN => gl_rom_n_1449);
  gl_rom_g34972 : ND4D0BWP7T port map(A1 => gl_rom_n_1334, A2 => gl_rom_n_1406, A3 => gl_rom_n_1416, A4 => gl_rom_n_1395, ZN => gl_rom_n_1448);
  gl_rom_g34973 : ND4D0BWP7T port map(A1 => gl_rom_n_1338, A2 => gl_rom_n_1339, A3 => gl_rom_n_1420, A4 => gl_rom_n_1332, ZN => gl_rom_n_1447);
  gl_rom_g34974 : AOI22D0BWP7T port map(A1 => gl_rom_n_1312, A2 => gl_rom_n_26, B1 => gl_rom_n_1314, B2 => gl_rom_n_27, ZN => gl_rom_n_1446);
  gl_rom_g34975 : AOI22D0BWP7T port map(A1 => gl_rom_n_1295, A2 => gl_rom_n_25, B1 => gl_rom_n_1297, B2 => gl_rom_n_28, ZN => gl_rom_n_1445);
  gl_rom_g34976 : AOI22D0BWP7T port map(A1 => gl_rom_n_1284, A2 => gl_rom_n_25, B1 => gl_rom_n_1290, B2 => gl_rom_n_28, ZN => gl_rom_n_1444);
  gl_rom_g34977 : AOI22D0BWP7T port map(A1 => gl_rom_n_1282, A2 => gl_rom_n_25, B1 => gl_rom_n_1285, B2 => gl_rom_n_28, ZN => gl_rom_n_1443);
  gl_rom_g34978 : AOI22D0BWP7T port map(A1 => gl_rom_n_1273, A2 => gl_rom_n_25, B1 => gl_rom_n_1276, B2 => gl_rom_n_28, ZN => gl_rom_n_1442);
  gl_rom_g34979 : AOI22D0BWP7T port map(A1 => gl_rom_n_1231, A2 => gl_rom_n_25, B1 => gl_rom_n_1264, B2 => gl_rom_n_28, ZN => gl_rom_n_1441);
  gl_rom_g34980 : AOI22D0BWP7T port map(A1 => gl_rom_n_1268, A2 => gl_rom_n_25, B1 => gl_rom_n_1270, B2 => gl_rom_n_28, ZN => gl_rom_n_1440);
  gl_rom_g34981 : AOI22D0BWP7T port map(A1 => gl_rom_n_1254, A2 => gl_rom_n_25, B1 => gl_rom_n_1255, B2 => gl_rom_n_28, ZN => gl_rom_n_1439);
  gl_rom_g34982 : AOI22D0BWP7T port map(A1 => gl_rom_n_1240, A2 => gl_rom_n_25, B1 => gl_rom_n_1244, B2 => gl_rom_n_28, ZN => gl_rom_n_1438);
  gl_rom_g34983 : AOI22D0BWP7T port map(A1 => gl_rom_n_1232, A2 => gl_rom_n_25, B1 => gl_rom_n_1233, B2 => gl_rom_n_28, ZN => gl_rom_n_1437);
  gl_rom_g34984 : AOI22D0BWP7T port map(A1 => gl_rom_n_1219, A2 => gl_rom_n_25, B1 => gl_rom_n_1222, B2 => gl_rom_n_28, ZN => gl_rom_n_1436);
  gl_rom_g34985 : AOI22D0BWP7T port map(A1 => gl_rom_n_1207, A2 => gl_rom_n_25, B1 => gl_rom_n_1212, B2 => gl_rom_n_28, ZN => gl_rom_n_1435);
  gl_rom_g34986 : AOI22D0BWP7T port map(A1 => gl_rom_n_1203, A2 => gl_rom_n_25, B1 => gl_rom_n_1205, B2 => gl_rom_n_28, ZN => gl_rom_n_1434);
  gl_rom_g34987 : AOI22D0BWP7T port map(A1 => gl_rom_n_1204, A2 => gl_rom_n_25, B1 => gl_rom_n_1206, B2 => gl_rom_n_28, ZN => gl_rom_n_1433);
  gl_rom_g34988 : AOI22D0BWP7T port map(A1 => gl_rom_n_1187, A2 => gl_rom_n_25, B1 => gl_rom_n_1189, B2 => gl_rom_n_28, ZN => gl_rom_n_1432);
  gl_rom_g34989 : AOI22D0BWP7T port map(A1 => gl_rom_n_1172, A2 => gl_rom_n_25, B1 => gl_rom_n_1180, B2 => gl_rom_n_28, ZN => gl_rom_n_1431);
  gl_rom_g34990 : AOI22D0BWP7T port map(A1 => gl_rom_n_1169, A2 => gl_rom_n_25, B1 => gl_rom_n_1173, B2 => gl_rom_n_28, ZN => gl_rom_n_1430);
  gl_rom_g34991 : AOI22D0BWP7T port map(A1 => gl_rom_n_1167, A2 => gl_rom_n_25, B1 => gl_rom_n_1168, B2 => gl_rom_n_28, ZN => gl_rom_n_1429);
  gl_rom_g34992 : AOI22D0BWP7T port map(A1 => gl_rom_n_1159, A2 => gl_rom_n_25, B1 => gl_rom_n_1160, B2 => gl_rom_n_28, ZN => gl_rom_n_1428);
  gl_rom_g34993 : AOI22D0BWP7T port map(A1 => gl_rom_n_1151, A2 => gl_rom_n_25, B1 => gl_rom_n_1165, B2 => gl_rom_n_28, ZN => gl_rom_n_1427);
  gl_rom_g34994 : AOI22D0BWP7T port map(A1 => gl_rom_n_1146, A2 => gl_rom_n_25, B1 => gl_rom_n_1149, B2 => gl_rom_n_28, ZN => gl_rom_n_1426);
  gl_rom_g34995 : AOI22D0BWP7T port map(A1 => gl_rom_n_1140, A2 => gl_rom_n_25, B1 => gl_rom_n_1142, B2 => gl_rom_n_28, ZN => gl_rom_n_1425);
  gl_rom_g34996 : AOI22D0BWP7T port map(A1 => gl_rom_n_1119, A2 => gl_rom_n_25, B1 => gl_rom_n_1120, B2 => gl_rom_n_28, ZN => gl_rom_n_1424);
  gl_rom_g34997 : AOI22D0BWP7T port map(A1 => gl_rom_n_1191, A2 => gl_rom_n_25, B1 => gl_rom_n_1085, B2 => gl_rom_n_28, ZN => gl_rom_n_1423);
  gl_rom_g34998 : AOI22D0BWP7T port map(A1 => gl_rom_n_1109, A2 => gl_rom_n_25, B1 => gl_rom_n_1115, B2 => gl_rom_n_28, ZN => gl_rom_n_1422);
  gl_rom_g34999 : AOI22D0BWP7T port map(A1 => gl_rom_n_1106, A2 => gl_rom_n_25, B1 => gl_rom_n_1110, B2 => gl_rom_n_28, ZN => gl_rom_n_1421);
  gl_rom_g35000 : AOI22D0BWP7T port map(A1 => gl_rom_n_1105, A2 => gl_rom_n_25, B1 => gl_rom_n_1107, B2 => gl_rom_n_28, ZN => gl_rom_n_1420);
  gl_rom_g35001 : AOI22D0BWP7T port map(A1 => gl_rom_n_1091, A2 => gl_rom_n_25, B1 => gl_rom_n_1093, B2 => gl_rom_n_28, ZN => gl_rom_n_1419);
  gl_rom_g35002 : AOI22D0BWP7T port map(A1 => gl_rom_n_1073, A2 => gl_rom_n_25, B1 => gl_rom_n_1075, B2 => gl_rom_n_28, ZN => gl_rom_n_1418);
  gl_rom_g35003 : AOI22D0BWP7T port map(A1 => gl_rom_n_1071, A2 => gl_rom_n_25, B1 => gl_rom_n_1072, B2 => gl_rom_n_28, ZN => gl_rom_n_1417);
  gl_rom_g35004 : AOI22D0BWP7T port map(A1 => gl_rom_n_1308, A2 => gl_rom_n_25, B1 => gl_rom_n_1067, B2 => gl_rom_n_28, ZN => gl_rom_n_1416);
  gl_rom_g35005 : AOI22D0BWP7T port map(A1 => gl_rom_n_1317, A2 => gl_rom_n_25, B1 => gl_rom_n_1190, B2 => gl_rom_n_28, ZN => gl_rom_n_1415);
  gl_rom_g35006 : AOI22D0BWP7T port map(A1 => gl_rom_n_1304, A2 => gl_rom_n_25, B1 => gl_rom_n_1307, B2 => gl_rom_n_28, ZN => gl_rom_n_1414);
  gl_rom_g35007 : AOI22D0BWP7T port map(A1 => gl_rom_n_1313, A2 => gl_rom_n_23, B1 => gl_rom_n_1315, B2 => gl_rom_n_30, ZN => gl_rom_n_1413);
  gl_rom_g35008 : AOI22D0BWP7T port map(A1 => gl_rom_n_1310, A2 => gl_rom_n_26, B1 => gl_rom_n_1311, B2 => gl_rom_n_27, ZN => gl_rom_n_1412);
  gl_rom_g35009 : AOI22D0BWP7T port map(A1 => gl_rom_n_1300, A2 => gl_rom_n_23, B1 => gl_rom_n_1306, B2 => gl_rom_n_30, ZN => gl_rom_n_1411);
  gl_rom_g35010 : AOI22D0BWP7T port map(A1 => gl_rom_n_1305, A2 => gl_rom_n_24, B1 => gl_rom_n_1309, B2 => gl_rom_n_29, ZN => gl_rom_n_1410);
  gl_rom_g35011 : AOI22D0BWP7T port map(A1 => gl_rom_n_1302, A2 => gl_rom_n_26, B1 => gl_rom_n_1303, B2 => gl_rom_n_27, ZN => gl_rom_n_1409);
  gl_rom_g35012 : AOI22D0BWP7T port map(A1 => gl_rom_n_1296, A2 => gl_rom_n_23, B1 => gl_rom_n_1299, B2 => gl_rom_n_30, ZN => gl_rom_n_1408);
  gl_rom_g35013 : AOI22D0BWP7T port map(A1 => gl_rom_n_1298, A2 => gl_rom_n_23, B1 => gl_rom_n_1301, B2 => gl_rom_n_30, ZN => gl_rom_n_1407);
  gl_rom_g35014 : AOI22D0BWP7T port map(A1 => gl_rom_n_1277, A2 => gl_rom_n_26, B1 => gl_rom_n_1291, B2 => gl_rom_n_27, ZN => gl_rom_n_1406);
  gl_rom_g35015 : AOI22D0BWP7T port map(A1 => gl_rom_n_1288, A2 => gl_rom_n_24, B1 => gl_rom_n_1292, B2 => gl_rom_n_29, ZN => gl_rom_n_1405);
  gl_rom_g35016 : AOI22D0BWP7T port map(A1 => gl_rom_n_1289, A2 => gl_rom_n_24, B1 => gl_rom_n_1293, B2 => gl_rom_n_29, ZN => gl_rom_n_1404);
  gl_rom_g35017 : AOI22D0BWP7T port map(A1 => gl_rom_n_1286, A2 => gl_rom_n_26, B1 => gl_rom_n_1287, B2 => gl_rom_n_27, ZN => gl_rom_n_1403);
  gl_rom_g35018 : AOI22D0BWP7T port map(A1 => gl_rom_n_1200, A2 => gl_rom_n_26, B1 => gl_rom_n_1262, B2 => gl_rom_n_27, ZN => gl_rom_n_1402);
  gl_rom_g35019 : AOI22D0BWP7T port map(A1 => gl_rom_n_1281, A2 => gl_rom_n_26, B1 => gl_rom_n_1283, B2 => gl_rom_n_27, ZN => gl_rom_n_1401);
  gl_rom_g35020 : AOI22D0BWP7T port map(A1 => gl_rom_n_1279, A2 => gl_rom_n_23, B1 => gl_rom_n_1280, B2 => gl_rom_n_30, ZN => gl_rom_n_1400);
  gl_rom_g35021 : AOI22D0BWP7T port map(A1 => gl_rom_n_1267, A2 => gl_rom_n_26, B1 => gl_rom_n_1275, B2 => gl_rom_n_27, ZN => gl_rom_n_1399);
  gl_rom_g35022 : AOI22D0BWP7T port map(A1 => gl_rom_n_1274, A2 => gl_rom_n_24, B1 => gl_rom_n_1278, B2 => gl_rom_n_29, ZN => gl_rom_n_1398);
  gl_rom_g35023 : AOI22D0BWP7T port map(A1 => gl_rom_n_1271, A2 => gl_rom_n_26, B1 => gl_rom_n_1272, B2 => gl_rom_n_27, ZN => gl_rom_n_1397);
  gl_rom_g35024 : AOI22D0BWP7T port map(A1 => gl_rom_n_1265, A2 => gl_rom_n_23, B1 => gl_rom_n_1269, B2 => gl_rom_n_30, ZN => gl_rom_n_1396);
  gl_rom_g35025 : AOI22D0BWP7T port map(A1 => gl_rom_n_1245, A2 => gl_rom_n_24, B1 => gl_rom_n_1261, B2 => gl_rom_n_29, ZN => gl_rom_n_1395);
  gl_rom_g35026 : AOI22D0BWP7T port map(A1 => gl_rom_n_1263, A2 => gl_rom_n_23, B1 => gl_rom_n_1266, B2 => gl_rom_n_30, ZN => gl_rom_n_1394);
  gl_rom_g35027 : AOI22D0BWP7T port map(A1 => gl_rom_n_1253, A2 => gl_rom_n_24, B1 => gl_rom_n_1259, B2 => gl_rom_n_29, ZN => gl_rom_n_1393);
  gl_rom_g35028 : AOI22D0BWP7T port map(A1 => gl_rom_n_1256, A2 => gl_rom_n_24, B1 => gl_rom_n_1258, B2 => gl_rom_n_29, ZN => gl_rom_n_1392);
  gl_rom_g35029 : AOI22D0BWP7T port map(A1 => gl_rom_n_1257, A2 => gl_rom_n_24, B1 => gl_rom_n_1260, B2 => gl_rom_n_29, ZN => gl_rom_n_1391);
  gl_rom_g35030 : AOI22D0BWP7T port map(A1 => gl_rom_n_1250, A2 => gl_rom_n_23, B1 => gl_rom_n_1252, B2 => gl_rom_n_30, ZN => gl_rom_n_1390);
  gl_rom_g35031 : AOI22D0BWP7T port map(A1 => gl_rom_n_1249, A2 => gl_rom_n_23, B1 => gl_rom_n_1251, B2 => gl_rom_n_30, ZN => gl_rom_n_1389);
  gl_rom_g35032 : AOI22D0BWP7T port map(A1 => gl_rom_n_1247, A2 => gl_rom_n_26, B1 => gl_rom_n_1248, B2 => gl_rom_n_27, ZN => gl_rom_n_1388);
  gl_rom_g35033 : AOI22D0BWP7T port map(A1 => gl_rom_n_1242, A2 => gl_rom_n_24, B1 => gl_rom_n_1246, B2 => gl_rom_n_29, ZN => gl_rom_n_1387);
  gl_rom_g35034 : AOI22D0BWP7T port map(A1 => gl_rom_n_1238, A2 => gl_rom_n_26, B1 => gl_rom_n_1243, B2 => gl_rom_n_27, ZN => gl_rom_n_1386);
  gl_rom_g35035 : AOI22D0BWP7T port map(A1 => gl_rom_n_1239, A2 => gl_rom_n_26, B1 => gl_rom_n_1241, B2 => gl_rom_n_27, ZN => gl_rom_n_1385);
  gl_rom_g35036 : AOI22D0BWP7T port map(A1 => gl_rom_n_1234, A2 => gl_rom_n_26, B1 => gl_rom_n_1236, B2 => gl_rom_n_27, ZN => gl_rom_n_1384);
  gl_rom_g35037 : AOI22D0BWP7T port map(A1 => gl_rom_n_1235, A2 => gl_rom_n_23, B1 => gl_rom_n_1237, B2 => gl_rom_n_30, ZN => gl_rom_n_1383);
  gl_rom_g35038 : AOI22D0BWP7T port map(A1 => gl_rom_n_1143, A2 => gl_rom_n_26, B1 => gl_rom_n_1148, B2 => gl_rom_n_27, ZN => gl_rom_n_1382);
  gl_rom_g35039 : AOI22D0BWP7T port map(A1 => gl_rom_n_1220, A2 => gl_rom_n_23, B1 => gl_rom_n_1227, B2 => gl_rom_n_30, ZN => gl_rom_n_1381);
  gl_rom_g35040 : AOI22D0BWP7T port map(A1 => gl_rom_n_1226, A2 => gl_rom_n_24, B1 => gl_rom_n_1229, B2 => gl_rom_n_29, ZN => gl_rom_n_1380);
  gl_rom_g35041 : AOI22D0BWP7T port map(A1 => gl_rom_n_1228, A2 => gl_rom_n_24, B1 => gl_rom_n_1230, B2 => gl_rom_n_29, ZN => gl_rom_n_1379);
  gl_rom_g35042 : AOI22D0BWP7T port map(A1 => gl_rom_n_1224, A2 => gl_rom_n_26, B1 => gl_rom_n_1225, B2 => gl_rom_n_27, ZN => gl_rom_n_1378);
  gl_rom_g35043 : AOI22D0BWP7T port map(A1 => gl_rom_n_1218, A2 => gl_rom_n_26, B1 => gl_rom_n_1221, B2 => gl_rom_n_27, ZN => gl_rom_n_1377);
  gl_rom_g35044 : AOI22D0BWP7T port map(A1 => gl_rom_n_1209, A2 => gl_rom_n_23, B1 => gl_rom_n_1213, B2 => gl_rom_n_30, ZN => gl_rom_n_1376);
  gl_rom_g35045 : AOI22D0BWP7T port map(A1 => gl_rom_n_1216, A2 => gl_rom_n_23, B1 => gl_rom_n_1217, B2 => gl_rom_n_30, ZN => gl_rom_n_1375);
  gl_rom_g35046 : AOI22D0BWP7T port map(A1 => gl_rom_n_1211, A2 => gl_rom_n_24, B1 => gl_rom_n_1215, B2 => gl_rom_n_29, ZN => gl_rom_n_1374);
  gl_rom_g35047 : AOI22D0BWP7T port map(A1 => gl_rom_n_1170, A2 => gl_rom_n_23, B1 => gl_rom_n_1199, B2 => gl_rom_n_30, ZN => gl_rom_n_1373);
  gl_rom_g35048 : AOI22D0BWP7T port map(A1 => gl_rom_n_1208, A2 => gl_rom_n_26, B1 => gl_rom_n_1210, B2 => gl_rom_n_27, ZN => gl_rom_n_1372);
  gl_rom_g35049 : AOI22D0BWP7T port map(A1 => gl_rom_n_1183, A2 => gl_rom_n_23, B1 => gl_rom_n_1197, B2 => gl_rom_n_30, ZN => gl_rom_n_1371);
  gl_rom_g35050 : AOI22D0BWP7T port map(A1 => gl_rom_n_1201, A2 => gl_rom_n_23, B1 => gl_rom_n_1202, B2 => gl_rom_n_30, ZN => gl_rom_n_1370);
  gl_rom_g35051 : AOI22D0BWP7T port map(A1 => gl_rom_n_1194, A2 => gl_rom_n_24, B1 => gl_rom_n_1198, B2 => gl_rom_n_29, ZN => gl_rom_n_1369);
  gl_rom_g35052 : AOI22D0BWP7T port map(A1 => gl_rom_n_1193, A2 => gl_rom_n_24, B1 => gl_rom_n_1196, B2 => gl_rom_n_29, ZN => gl_rom_n_1368);
  gl_rom_g35053 : AOI22D0BWP7T port map(A1 => gl_rom_n_1318, A2 => gl_rom_n_23, B1 => gl_rom_n_1192, B2 => gl_rom_n_30, ZN => gl_rom_n_1367);
  gl_rom_g35054 : AOI22D0BWP7T port map(A1 => gl_rom_n_1063, A2 => gl_rom_n_24, B1 => gl_rom_n_1195, B2 => gl_rom_n_29, ZN => gl_rom_n_1366);
  gl_rom_g35055 : AOI22D0BWP7T port map(A1 => gl_rom_n_1185, A2 => gl_rom_n_26, B1 => gl_rom_n_1188, B2 => gl_rom_n_27, ZN => gl_rom_n_1365);
  gl_rom_g35056 : AOI22D0BWP7T port map(A1 => gl_rom_n_1184, A2 => gl_rom_n_26, B1 => gl_rom_n_1186, B2 => gl_rom_n_27, ZN => gl_rom_n_1364);
  gl_rom_g35057 : AOI22D0BWP7T port map(A1 => gl_rom_n_1177, A2 => gl_rom_n_23, B1 => gl_rom_n_1181, B2 => gl_rom_n_30, ZN => gl_rom_n_1363);
  gl_rom_g35058 : AOI22D0BWP7T port map(A1 => gl_rom_n_1179, A2 => gl_rom_n_24, B1 => gl_rom_n_1182, B2 => gl_rom_n_29, ZN => gl_rom_n_1362);
  gl_rom_g35059 : AOI22D0BWP7T port map(A1 => gl_rom_n_1087, A2 => gl_rom_n_23, B1 => gl_rom_n_1178, B2 => gl_rom_n_30, ZN => gl_rom_n_1361);
  gl_rom_g35060 : AOI22D0BWP7T port map(A1 => gl_rom_n_1175, A2 => gl_rom_n_26, B1 => gl_rom_n_1176, B2 => gl_rom_n_27, ZN => gl_rom_n_1360);
  gl_rom_g35061 : AOI22D0BWP7T port map(A1 => gl_rom_n_1171, A2 => gl_rom_n_23, B1 => gl_rom_n_1174, B2 => gl_rom_n_30, ZN => gl_rom_n_1359);
  gl_rom_g35062 : AOI22D0BWP7T port map(A1 => gl_rom_n_1156, A2 => gl_rom_n_23, B1 => gl_rom_n_1163, B2 => gl_rom_n_30, ZN => gl_rom_n_1358);
  gl_rom_g35063 : AOI22D0BWP7T port map(A1 => gl_rom_n_1161, A2 => gl_rom_n_24, B1 => gl_rom_n_1164, B2 => gl_rom_n_29, ZN => gl_rom_n_1357);
  gl_rom_g35064 : AOI22D0BWP7T port map(A1 => gl_rom_n_1162, A2 => gl_rom_n_24, B1 => gl_rom_n_1166, B2 => gl_rom_n_29, ZN => gl_rom_n_1356);
  gl_rom_g35065 : AOI22D0BWP7T port map(A1 => gl_rom_n_1153, A2 => gl_rom_n_26, B1 => gl_rom_n_1157, B2 => gl_rom_n_27, ZN => gl_rom_n_1355);
  gl_rom_g35066 : AOI22D0BWP7T port map(A1 => gl_rom_n_1155, A2 => gl_rom_n_23, B1 => gl_rom_n_1158, B2 => gl_rom_n_30, ZN => gl_rom_n_1354);
  gl_rom_g35067 : AOI22D0BWP7T port map(A1 => gl_rom_n_1108, A2 => gl_rom_n_24, B1 => gl_rom_n_1139, B2 => gl_rom_n_29, ZN => gl_rom_n_1353);
  gl_rom_g35068 : AOI22D0BWP7T port map(A1 => gl_rom_n_1152, A2 => gl_rom_n_26, B1 => gl_rom_n_1154, B2 => gl_rom_n_27, ZN => gl_rom_n_1352);
  gl_rom_g35069 : AOI22D0BWP7T port map(A1 => gl_rom_n_1118, A2 => gl_rom_n_24, B1 => gl_rom_n_1135, B2 => gl_rom_n_29, ZN => gl_rom_n_1351);
  gl_rom_g35070 : AOI22D0BWP7T port map(A1 => gl_rom_n_1214, A2 => gl_rom_n_26, B1 => gl_rom_n_1223, B2 => gl_rom_n_27, ZN => gl_rom_n_1350);
  gl_rom_g35071 : AOI22D0BWP7T port map(A1 => gl_rom_n_1147, A2 => gl_rom_n_24, B1 => gl_rom_n_1150, B2 => gl_rom_n_29, ZN => gl_rom_n_1349);
  gl_rom_g35072 : AOI22D0BWP7T port map(A1 => gl_rom_n_1144, A2 => gl_rom_n_26, B1 => gl_rom_n_1145, B2 => gl_rom_n_27, ZN => gl_rom_n_1348);
  gl_rom_g35073 : AOI22D0BWP7T port map(A1 => gl_rom_n_1138, A2 => gl_rom_n_23, B1 => gl_rom_n_1141, B2 => gl_rom_n_30, ZN => gl_rom_n_1347);
  gl_rom_g35074 : AOI22D0BWP7T port map(A1 => gl_rom_n_1136, A2 => gl_rom_n_23, B1 => gl_rom_n_1137, B2 => gl_rom_n_30, ZN => gl_rom_n_1346);
  gl_rom_g35075 : AOI22D0BWP7T port map(A1 => gl_rom_n_1128, A2 => gl_rom_n_24, B1 => gl_rom_n_1131, B2 => gl_rom_n_29, ZN => gl_rom_n_1345);
  gl_rom_g35076 : AOI22D0BWP7T port map(A1 => gl_rom_n_1129, A2 => gl_rom_n_24, B1 => gl_rom_n_1132, B2 => gl_rom_n_29, ZN => gl_rom_n_1344);
  gl_rom_g35077 : AOI22D0BWP7T port map(A1 => gl_rom_n_1130, A2 => gl_rom_n_24, B1 => gl_rom_n_1134, B2 => gl_rom_n_29, ZN => gl_rom_n_1343);
  gl_rom_g35078 : AOI22D0BWP7T port map(A1 => gl_rom_n_1126, A2 => gl_rom_n_26, B1 => gl_rom_n_1127, B2 => gl_rom_n_27, ZN => gl_rom_n_1342);
  gl_rom_g35079 : AOI22D0BWP7T port map(A1 => gl_rom_n_1125, A2 => gl_rom_n_24, B1 => gl_rom_n_1133, B2 => gl_rom_n_29, ZN => gl_rom_n_1341);
  gl_rom_g35080 : AOI22D0BWP7T port map(A1 => gl_rom_n_1122, A2 => gl_rom_n_23, B1 => gl_rom_n_1124, B2 => gl_rom_n_30, ZN => gl_rom_n_1340);
  gl_rom_g35081 : AOI22D0BWP7T port map(A1 => gl_rom_n_1121, A2 => gl_rom_n_26, B1 => gl_rom_n_1123, B2 => gl_rom_n_27, ZN => gl_rom_n_1339);
  gl_rom_g35082 : AOI22D0BWP7T port map(A1 => gl_rom_n_1113, A2 => gl_rom_n_23, B1 => gl_rom_n_1116, B2 => gl_rom_n_30, ZN => gl_rom_n_1338);
  gl_rom_g35083 : AOI22D0BWP7T port map(A1 => gl_rom_n_1114, A2 => gl_rom_n_24, B1 => gl_rom_n_1117, B2 => gl_rom_n_29, ZN => gl_rom_n_1337);
  gl_rom_g35084 : AOI22D0BWP7T port map(A1 => gl_rom_n_1111, A2 => gl_rom_n_23, B1 => gl_rom_n_1112, B2 => gl_rom_n_30, ZN => gl_rom_n_1336);
  gl_rom_g35085 : AOI22D0BWP7T port map(A1 => gl_rom_n_1103, A2 => gl_rom_n_26, B1 => gl_rom_n_1104, B2 => gl_rom_n_27, ZN => gl_rom_n_1335);
  gl_rom_g35086 : AOI22D0BWP7T port map(A1 => gl_rom_n_1084, A2 => gl_rom_n_23, B1 => gl_rom_n_1099, B2 => gl_rom_n_30, ZN => gl_rom_n_1334);
  gl_rom_g35087 : AOI22D0BWP7T port map(A1 => gl_rom_n_1094, A2 => gl_rom_n_23, B1 => gl_rom_n_1101, B2 => gl_rom_n_30, ZN => gl_rom_n_1333);
  gl_rom_g35088 : AOI22D0BWP7T port map(A1 => gl_rom_n_1096, A2 => gl_rom_n_24, B1 => gl_rom_n_1100, B2 => gl_rom_n_29, ZN => gl_rom_n_1332);
  gl_rom_g35089 : AOI22D0BWP7T port map(A1 => gl_rom_n_1098, A2 => gl_rom_n_24, B1 => gl_rom_n_1102, B2 => gl_rom_n_29, ZN => gl_rom_n_1331);
  gl_rom_g35090 : AOI22D0BWP7T port map(A1 => gl_rom_n_1095, A2 => gl_rom_n_26, B1 => gl_rom_n_1097, B2 => gl_rom_n_27, ZN => gl_rom_n_1330);
  gl_rom_g35091 : AOI22D0BWP7T port map(A1 => gl_rom_n_1090, A2 => gl_rom_n_26, B1 => gl_rom_n_1092, B2 => gl_rom_n_27, ZN => gl_rom_n_1329);
  gl_rom_g35092 : AOI22D0BWP7T port map(A1 => gl_rom_n_1076, A2 => gl_rom_n_26, B1 => gl_rom_n_1083, B2 => gl_rom_n_27, ZN => gl_rom_n_1328);
  gl_rom_g35093 : AOI22D0BWP7T port map(A1 => gl_rom_n_1088, A2 => gl_rom_n_23, B1 => gl_rom_n_1089, B2 => gl_rom_n_30, ZN => gl_rom_n_1327);
  gl_rom_g35094 : AOI22D0BWP7T port map(A1 => gl_rom_n_1080, A2 => gl_rom_n_23, B1 => gl_rom_n_1082, B2 => gl_rom_n_30, ZN => gl_rom_n_1326);
  gl_rom_g35095 : AOI22D0BWP7T port map(A1 => gl_rom_n_1081, A2 => gl_rom_n_24, B1 => gl_rom_n_1086, B2 => gl_rom_n_29, ZN => gl_rom_n_1325);
  gl_rom_g35096 : AOI22D0BWP7T port map(A1 => gl_rom_n_1078, A2 => gl_rom_n_26, B1 => gl_rom_n_1079, B2 => gl_rom_n_27, ZN => gl_rom_n_1324);
  gl_rom_g35097 : AOI22D0BWP7T port map(A1 => gl_rom_n_1074, A2 => gl_rom_n_23, B1 => gl_rom_n_1077, B2 => gl_rom_n_30, ZN => gl_rom_n_1323);
  gl_rom_g35098 : AOI22D0BWP7T port map(A1 => gl_rom_n_1294, A2 => gl_rom_n_26, B1 => gl_rom_n_1065, B2 => gl_rom_n_27, ZN => gl_rom_n_1322);
  gl_rom_g35099 : AOI22D0BWP7T port map(A1 => gl_rom_n_1316, A2 => gl_rom_n_24, B1 => gl_rom_n_1069, B2 => gl_rom_n_29, ZN => gl_rom_n_1321);
  gl_rom_g35100 : AOI22D0BWP7T port map(A1 => gl_rom_n_1064, A2 => gl_rom_n_24, B1 => gl_rom_n_1068, B2 => gl_rom_n_29, ZN => gl_rom_n_1320);
  gl_rom_g35101 : AOI22D0BWP7T port map(A1 => gl_rom_n_1066, A2 => gl_rom_n_24, B1 => gl_rom_n_1070, B2 => gl_rom_n_29, ZN => gl_rom_n_1319);
  gl_rom_g35102 : ND4D0BWP7T port map(A1 => gl_rom_n_546, A2 => gl_rom_n_294, A3 => gl_rom_n_549, A4 => gl_rom_n_547, ZN => gl_rom_n_1318);
  gl_rom_g35103 : ND4D0BWP7T port map(A1 => gl_rom_n_1056, A2 => gl_rom_n_1060, A3 => gl_rom_n_1059, A4 => gl_rom_n_1057, ZN => gl_rom_n_1317);
  gl_rom_g35104 : ND4D0BWP7T port map(A1 => gl_rom_n_1052, A2 => gl_rom_n_1036, A3 => gl_rom_n_1046, A4 => gl_rom_n_1033, ZN => gl_rom_n_1316);
  gl_rom_g35105 : ND4D0BWP7T port map(A1 => gl_rom_n_1047, A2 => gl_rom_n_1051, A3 => gl_rom_n_1050, A4 => gl_rom_n_1048, ZN => gl_rom_n_1315);
  gl_rom_g35106 : ND4D0BWP7T port map(A1 => gl_rom_n_1049, A2 => gl_rom_n_1041, A3 => gl_rom_n_1045, A4 => gl_rom_n_1039, ZN => gl_rom_n_1314);
  gl_rom_g35107 : ND4D0BWP7T port map(A1 => gl_rom_n_1043, A2 => gl_rom_n_1044, A3 => gl_rom_n_1040, A4 => gl_rom_n_1038, ZN => gl_rom_n_1313);
  gl_rom_g35108 : ND4D0BWP7T port map(A1 => gl_rom_n_1030, A2 => gl_rom_n_1034, A3 => gl_rom_n_1026, A4 => gl_rom_n_1025, ZN => gl_rom_n_1312);
  gl_rom_g35109 : ND4D0BWP7T port map(A1 => gl_rom_n_1032, A2 => gl_rom_n_1035, A3 => gl_rom_n_1037, A4 => gl_rom_n_1031, ZN => gl_rom_n_1311);
  gl_rom_g35110 : ND4D0BWP7T port map(A1 => gl_rom_n_1024, A2 => gl_rom_n_1027, A3 => gl_rom_n_1029, A4 => gl_rom_n_1023, ZN => gl_rom_n_1310);
  gl_rom_g35111 : ND4D0BWP7T port map(A1 => gl_rom_n_1018, A2 => gl_rom_n_1020, A3 => gl_rom_n_1022, A4 => gl_rom_n_1016, ZN => gl_rom_n_1309);
  gl_rom_g35112 : ND4D0BWP7T port map(A1 => gl_rom_n_990, A2 => gl_rom_n_1010, A3 => gl_rom_n_1017, A4 => gl_rom_n_982, ZN => gl_rom_n_1308);
  gl_rom_g35113 : ND4D0BWP7T port map(A1 => gl_rom_n_1019, A2 => gl_rom_n_1012, A3 => gl_rom_n_1015, A4 => gl_rom_n_1007, ZN => gl_rom_n_1307);
  gl_rom_g35114 : ND4D0BWP7T port map(A1 => gl_rom_n_1005, A2 => gl_rom_n_1014, A3 => gl_rom_n_1004, A4 => gl_rom_n_998, ZN => gl_rom_n_1306);
  gl_rom_g35115 : ND4D0BWP7T port map(A1 => gl_rom_n_1009, A2 => gl_rom_n_1011, A3 => gl_rom_n_1013, A4 => gl_rom_n_1008, ZN => gl_rom_n_1305);
  gl_rom_g35116 : ND4D0BWP7T port map(A1 => gl_rom_n_1002, A2 => gl_rom_n_996, A3 => gl_rom_n_1000, A4 => gl_rom_n_993, ZN => gl_rom_n_1304);
  gl_rom_g35117 : ND4D0BWP7T port map(A1 => gl_rom_n_999, A2 => gl_rom_n_1006, A3 => gl_rom_n_1003, A4 => gl_rom_n_1001, ZN => gl_rom_n_1303);
  gl_rom_g35118 : ND4D0BWP7T port map(A1 => gl_rom_n_992, A2 => gl_rom_n_997, A3 => gl_rom_n_995, A4 => gl_rom_n_994, ZN => gl_rom_n_1302);
  gl_rom_g35119 : ND4D0BWP7T port map(A1 => gl_rom_n_986, A2 => gl_rom_n_989, A3 => gl_rom_n_991, A4 => gl_rom_n_984, ZN => gl_rom_n_1301);
  gl_rom_g35120 : ND4D0BWP7T port map(A1 => gl_rom_n_970, A2 => gl_rom_n_985, A3 => gl_rom_n_975, A4 => gl_rom_n_965, ZN => gl_rom_n_1300);
  gl_rom_g35121 : ND4D0BWP7T port map(A1 => gl_rom_n_987, A2 => gl_rom_n_979, A3 => gl_rom_n_983, A4 => gl_rom_n_977, ZN => gl_rom_n_1299);
  gl_rom_g35122 : ND4D0BWP7T port map(A1 => gl_rom_n_980, A2 => gl_rom_n_981, A3 => gl_rom_n_978, A4 => gl_rom_n_976, ZN => gl_rom_n_1298);
  gl_rom_g35123 : ND4D0BWP7T port map(A1 => gl_rom_n_967, A2 => gl_rom_n_974, A3 => gl_rom_n_972, A4 => gl_rom_n_969, ZN => gl_rom_n_1297);
  gl_rom_g35124 : ND4D0BWP7T port map(A1 => gl_rom_n_971, A2 => gl_rom_n_964, A3 => gl_rom_n_968, A4 => gl_rom_n_962, ZN => gl_rom_n_1296);
  gl_rom_g35125 : ND4D0BWP7T port map(A1 => gl_rom_n_963, A2 => gl_rom_n_960, A3 => gl_rom_n_966, A4 => gl_rom_n_961, ZN => gl_rom_n_1295);
  gl_rom_g35126 : ND4D0BWP7T port map(A1 => gl_rom_n_952, A2 => gl_rom_n_902, A3 => gl_rom_n_925, A4 => gl_rom_n_865, ZN => gl_rom_n_1294);
  gl_rom_g35127 : ND4D0BWP7T port map(A1 => gl_rom_n_956, A2 => gl_rom_n_959, A3 => gl_rom_n_958, A4 => gl_rom_n_955, ZN => gl_rom_n_1293);
  gl_rom_g35128 : ND4D0BWP7T port map(A1 => gl_rom_n_946, A2 => gl_rom_n_957, A3 => gl_rom_n_954, A4 => gl_rom_n_949, ZN => gl_rom_n_1292);
  gl_rom_g35129 : ND4D0BWP7T port map(A1 => gl_rom_n_950, A2 => gl_rom_n_928, A3 => gl_rom_n_943, A4 => gl_rom_n_910, ZN => gl_rom_n_1291);
  gl_rom_g35130 : ND4D0BWP7T port map(A1 => gl_rom_n_933, A2 => gl_rom_n_953, A3 => gl_rom_n_947, A4 => gl_rom_n_939, ZN => gl_rom_n_1290);
  gl_rom_g35131 : ND4D0BWP7T port map(A1 => gl_rom_n_948, A2 => gl_rom_n_951, A3 => gl_rom_n_945, A4 => gl_rom_n_944, ZN => gl_rom_n_1289);
  gl_rom_g35132 : ND4D0BWP7T port map(A1 => gl_rom_n_941, A2 => gl_rom_n_935, A3 => gl_rom_n_936, A4 => gl_rom_n_931, ZN => gl_rom_n_1288);
  gl_rom_g35133 : ND4D0BWP7T port map(A1 => gl_rom_n_938, A2 => gl_rom_n_940, A3 => gl_rom_n_942, A4 => gl_rom_n_937, ZN => gl_rom_n_1287);
  gl_rom_g35134 : ND4D0BWP7T port map(A1 => gl_rom_n_930, A2 => gl_rom_n_932, A3 => gl_rom_n_934, A4 => gl_rom_n_929, ZN => gl_rom_n_1286);
  gl_rom_g35135 : ND4D0BWP7T port map(A1 => gl_rom_n_927, A2 => gl_rom_n_923, A3 => gl_rom_n_926, A4 => gl_rom_n_922, ZN => gl_rom_n_1285);
  gl_rom_g35136 : ND4D0BWP7T port map(A1 => gl_rom_n_917, A2 => gl_rom_n_901, A3 => gl_rom_n_919, A4 => gl_rom_n_909, ZN => gl_rom_n_1284);
  gl_rom_g35137 : ND4D0BWP7T port map(A1 => gl_rom_n_916, A2 => gl_rom_n_921, A3 => gl_rom_n_924, A4 => gl_rom_n_915, ZN => gl_rom_n_1283);
  gl_rom_g35138 : ND4D0BWP7T port map(A1 => gl_rom_n_914, A2 => gl_rom_n_918, A3 => gl_rom_n_920, A4 => gl_rom_n_913, ZN => gl_rom_n_1282);
  gl_rom_g35139 : ND4D0BWP7T port map(A1 => gl_rom_n_906, A2 => gl_rom_n_898, A3 => gl_rom_n_907, A4 => gl_rom_n_900, ZN => gl_rom_n_1281);
  gl_rom_g35140 : ND4D0BWP7T port map(A1 => gl_rom_n_908, A2 => gl_rom_n_904, A3 => gl_rom_n_912, A4 => gl_rom_n_905, ZN => gl_rom_n_1280);
  gl_rom_g35141 : ND4D0BWP7T port map(A1 => gl_rom_n_897, A2 => gl_rom_n_899, A3 => gl_rom_n_903, A4 => gl_rom_n_896, ZN => gl_rom_n_1279);
  gl_rom_g35142 : ND4D0BWP7T port map(A1 => gl_rom_n_891, A2 => gl_rom_n_894, A3 => gl_rom_n_895, A4 => gl_rom_n_889, ZN => gl_rom_n_1278);
  gl_rom_g35143 : ND4D0BWP7T port map(A1 => gl_rom_n_879, A2 => gl_rom_n_846, A3 => gl_rom_n_893, A4 => gl_rom_n_864, ZN => gl_rom_n_1277);
  gl_rom_g35144 : ND4D0BWP7T port map(A1 => gl_rom_n_892, A2 => gl_rom_n_885, A3 => gl_rom_n_890, A4 => gl_rom_n_880, ZN => gl_rom_n_1276);
  gl_rom_g35145 : ND4D0BWP7T port map(A1 => gl_rom_n_872, A2 => gl_rom_n_888, A3 => gl_rom_n_887, A4 => gl_rom_n_876, ZN => gl_rom_n_1275);
  gl_rom_g35146 : ND4D0BWP7T port map(A1 => gl_rom_n_884, A2 => gl_rom_n_886, A3 => gl_rom_n_883, A4 => gl_rom_n_882, ZN => gl_rom_n_1274);
  gl_rom_g35147 : ND4D0BWP7T port map(A1 => gl_rom_n_878, A2 => gl_rom_n_871, A3 => gl_rom_n_874, A4 => gl_rom_n_867, ZN => gl_rom_n_1273);
  gl_rom_g35148 : ND4D0BWP7T port map(A1 => gl_rom_n_873, A2 => gl_rom_n_881, A3 => gl_rom_n_877, A4 => gl_rom_n_875, ZN => gl_rom_n_1272);
  gl_rom_g35149 : ND4D0BWP7T port map(A1 => gl_rom_n_869, A2 => gl_rom_n_870, A3 => gl_rom_n_868, A4 => gl_rom_n_866, ZN => gl_rom_n_1271);
  gl_rom_g35150 : ND4D0BWP7T port map(A1 => gl_rom_n_857, A2 => gl_rom_n_860, A3 => gl_rom_n_863, A4 => gl_rom_n_855, ZN => gl_rom_n_1270);
  gl_rom_g35151 : ND4D0BWP7T port map(A1 => gl_rom_n_859, A2 => gl_rom_n_853, A3 => gl_rom_n_856, A4 => gl_rom_n_848, ZN => gl_rom_n_1269);
  gl_rom_g35152 : ND4D0BWP7T port map(A1 => gl_rom_n_850, A2 => gl_rom_n_852, A3 => gl_rom_n_854, A4 => gl_rom_n_849, ZN => gl_rom_n_1268);
  gl_rom_g35153 : ND4D0BWP7T port map(A1 => gl_rom_n_851, A2 => gl_rom_n_838, A3 => gl_rom_n_858, A4 => gl_rom_n_845, ZN => gl_rom_n_1267);
  gl_rom_g35154 : ND4D0BWP7T port map(A1 => gl_rom_n_841, A2 => gl_rom_n_843, A3 => gl_rom_n_847, A4 => gl_rom_n_840, ZN => gl_rom_n_1266);
  gl_rom_g35155 : ND4D0BWP7T port map(A1 => gl_rom_n_837, A2 => gl_rom_n_842, A3 => gl_rom_n_844, A4 => gl_rom_n_835, ZN => gl_rom_n_1265);
  gl_rom_g35156 : ND4D0BWP7T port map(A1 => gl_rom_n_798, A2 => gl_rom_n_742, A3 => gl_rom_n_824, A4 => gl_rom_n_768, ZN => gl_rom_n_1264);
  gl_rom_g35157 : ND4D0BWP7T port map(A1 => gl_rom_n_834, A2 => gl_rom_n_836, A3 => gl_rom_n_839, A4 => gl_rom_n_833, ZN => gl_rom_n_1263);
  gl_rom_g35158 : ND4D0BWP7T port map(A1 => gl_rom_n_816, A2 => gl_rom_n_861, A3 => gl_rom_n_743, A4 => gl_rom_n_706, ZN => gl_rom_n_1262);
  gl_rom_g35159 : ND4D0BWP7T port map(A1 => gl_rom_n_811, A2 => gl_rom_n_783, A3 => gl_rom_n_829, A4 => gl_rom_n_800, ZN => gl_rom_n_1261);
  gl_rom_g35160 : ND4D0BWP7T port map(A1 => gl_rom_n_828, A2 => gl_rom_n_831, A3 => gl_rom_n_832, A4 => gl_rom_n_826, ZN => gl_rom_n_1260);
  gl_rom_g35161 : ND4D0BWP7T port map(A1 => gl_rom_n_817, A2 => gl_rom_n_827, A3 => gl_rom_n_814, A4 => gl_rom_n_1062, ZN => gl_rom_n_1259);
  gl_rom_g35162 : ND4D0BWP7T port map(A1 => gl_rom_n_825, A2 => gl_rom_n_820, A3 => gl_rom_n_830, A4 => gl_rom_n_822, ZN => gl_rom_n_1258);
  gl_rom_g35163 : ND4D0BWP7T port map(A1 => gl_rom_n_819, A2 => gl_rom_n_823, A3 => gl_rom_n_821, A4 => gl_rom_n_818, ZN => gl_rom_n_1257);
  gl_rom_g35164 : ND4D0BWP7T port map(A1 => gl_rom_n_815, A2 => gl_rom_n_807, A3 => gl_rom_n_810, A4 => gl_rom_n_803, ZN => gl_rom_n_1256);
  gl_rom_g35165 : ND4D0BWP7T port map(A1 => gl_rom_n_812, A2 => gl_rom_n_813, A3 => gl_rom_n_809, A4 => gl_rom_n_808, ZN => gl_rom_n_1255);
  gl_rom_g35166 : ND4D0BWP7T port map(A1 => gl_rom_n_802, A2 => gl_rom_n_805, A3 => gl_rom_n_804, A4 => gl_rom_n_801, ZN => gl_rom_n_1254);
  gl_rom_g35167 : ND4D0BWP7T port map(A1 => gl_rom_n_791, A2 => gl_rom_n_797, A3 => gl_rom_n_782, A4 => gl_rom_n_779, ZN => gl_rom_n_1253);
  gl_rom_g35168 : ND4D0BWP7T port map(A1 => gl_rom_n_799, A2 => gl_rom_n_794, A3 => gl_rom_n_796, A4 => gl_rom_n_793, ZN => gl_rom_n_1252);
  gl_rom_g35169 : ND4D0BWP7T port map(A1 => gl_rom_n_785, A2 => gl_rom_n_795, A3 => gl_rom_n_792, A4 => gl_rom_n_788, ZN => gl_rom_n_1251);
  gl_rom_g35170 : ND4D0BWP7T port map(A1 => gl_rom_n_787, A2 => gl_rom_n_789, A3 => gl_rom_n_790, A4 => gl_rom_n_786, ZN => gl_rom_n_1250);
  gl_rom_g35171 : ND4D0BWP7T port map(A1 => gl_rom_n_770, A2 => gl_rom_n_781, A3 => gl_rom_n_777, A4 => gl_rom_n_774, ZN => gl_rom_n_1249);
  gl_rom_g35172 : ND4D0BWP7T port map(A1 => gl_rom_n_784, A2 => gl_rom_n_778, A3 => gl_rom_n_780, A4 => gl_rom_n_776, ZN => gl_rom_n_1248);
  gl_rom_g35173 : ND4D0BWP7T port map(A1 => gl_rom_n_771, A2 => gl_rom_n_775, A3 => gl_rom_n_773, A4 => gl_rom_n_769, ZN => gl_rom_n_1247);
  gl_rom_g35174 : ND4D0BWP7T port map(A1 => gl_rom_n_765, A2 => gl_rom_n_766, A3 => gl_rom_n_763, A4 => gl_rom_n_762, ZN => gl_rom_n_1246);
  gl_rom_g35175 : ND4D0BWP7T port map(A1 => gl_rom_n_752, A2 => gl_rom_n_726, A3 => gl_rom_n_767, A4 => gl_rom_n_735, ZN => gl_rom_n_1245);
  gl_rom_g35176 : ND4D0BWP7T port map(A1 => gl_rom_n_761, A2 => gl_rom_n_764, A3 => gl_rom_n_758, A4 => gl_rom_n_754, ZN => gl_rom_n_1244);
  gl_rom_g35177 : ND4D0BWP7T port map(A1 => gl_rom_n_744, A2 => gl_rom_n_751, A3 => gl_rom_n_760, A4 => gl_rom_n_732, ZN => gl_rom_n_1243);
  gl_rom_g35178 : ND4D0BWP7T port map(A1 => gl_rom_n_755, A2 => gl_rom_n_759, A3 => gl_rom_n_757, A4 => gl_rom_n_753, ZN => gl_rom_n_1242);
  gl_rom_g35179 : ND4D0BWP7T port map(A1 => gl_rom_n_750, A2 => gl_rom_n_746, A3 => gl_rom_n_748, A4 => gl_rom_n_745, ZN => gl_rom_n_1241);
  gl_rom_g35180 : ND4D0BWP7T port map(A1 => gl_rom_n_740, A2 => gl_rom_n_747, A3 => gl_rom_n_749, A4 => gl_rom_n_736, ZN => gl_rom_n_1240);
  gl_rom_g35181 : ND4D0BWP7T port map(A1 => gl_rom_n_739, A2 => gl_rom_n_741, A3 => gl_rom_n_738, A4 => gl_rom_n_737, ZN => gl_rom_n_1239);
  gl_rom_g35182 : ND4D0BWP7T port map(A1 => gl_rom_n_708, A2 => gl_rom_n_727, A3 => gl_rom_n_722, A4 => gl_rom_n_712, ZN => gl_rom_n_1238);
  gl_rom_g35183 : ND4D0BWP7T port map(A1 => gl_rom_n_733, A2 => gl_rom_n_734, A3 => gl_rom_n_730, A4 => gl_rom_n_728, ZN => gl_rom_n_1237);
  gl_rom_g35184 : ND4D0BWP7T port map(A1 => gl_rom_n_724, A2 => gl_rom_n_729, A3 => gl_rom_n_731, A4 => gl_rom_n_719, ZN => gl_rom_n_1236);
  gl_rom_g35185 : ND4D0BWP7T port map(A1 => gl_rom_n_721, A2 => gl_rom_n_723, A3 => gl_rom_n_725, A4 => gl_rom_n_720, ZN => gl_rom_n_1235);
  gl_rom_g35186 : ND4D0BWP7T port map(A1 => gl_rom_n_705, A2 => gl_rom_n_716, A3 => gl_rom_n_714, A4 => gl_rom_n_710, ZN => gl_rom_n_1234);
  gl_rom_g35187 : ND4D0BWP7T port map(A1 => gl_rom_n_715, A2 => gl_rom_n_718, A3 => gl_rom_n_717, A4 => gl_rom_n_713, ZN => gl_rom_n_1233);
  gl_rom_g35188 : ND4D0BWP7T port map(A1 => gl_rom_n_709, A2 => gl_rom_n_711, A3 => gl_rom_n_707, A4 => gl_rom_n_704, ZN => gl_rom_n_1232);
  gl_rom_g35189 : ND4D0BWP7T port map(A1 => gl_rom_n_703, A2 => gl_rom_n_639, A3 => gl_rom_n_698, A4 => gl_rom_n_636, ZN => gl_rom_n_1231);
  gl_rom_g35190 : ND4D0BWP7T port map(A1 => gl_rom_n_699, A2 => gl_rom_n_702, A3 => gl_rom_n_701, A4 => gl_rom_n_696, ZN => gl_rom_n_1230);
  gl_rom_g35191 : ND4D0BWP7T port map(A1 => gl_rom_n_688, A2 => gl_rom_n_700, A3 => gl_rom_n_697, A4 => gl_rom_n_691, ZN => gl_rom_n_1229);
  gl_rom_g35192 : ND4D0BWP7T port map(A1 => gl_rom_n_690, A2 => gl_rom_n_692, A3 => gl_rom_n_694, A4 => gl_rom_n_687, ZN => gl_rom_n_1228);
  gl_rom_g35193 : ND4D0BWP7T port map(A1 => gl_rom_n_695, A2 => gl_rom_n_683, A3 => gl_rom_n_689, A4 => gl_rom_n_672, ZN => gl_rom_n_1227);
  gl_rom_g35194 : ND4D0BWP7T port map(A1 => gl_rom_n_675, A2 => gl_rom_n_686, A3 => gl_rom_n_682, A4 => gl_rom_n_678, ZN => gl_rom_n_1226);
  gl_rom_g35195 : ND4D0BWP7T port map(A1 => gl_rom_n_680, A2 => gl_rom_n_685, A3 => gl_rom_n_684, A4 => gl_rom_n_681, ZN => gl_rom_n_1225);
  gl_rom_g35196 : ND4D0BWP7T port map(A1 => gl_rom_n_676, A2 => gl_rom_n_673, A3 => gl_rom_n_677, A4 => gl_rom_n_674, ZN => gl_rom_n_1224);
  gl_rom_g35197 : ND4D0BWP7T port map(A1 => gl_rom_n_693, A2 => gl_rom_n_669, A3 => gl_rom_n_679, A4 => gl_rom_n_652, ZN => gl_rom_n_1223);
  gl_rom_g35198 : ND4D0BWP7T port map(A1 => gl_rom_n_666, A2 => gl_rom_n_671, A3 => gl_rom_n_670, A4 => gl_rom_n_667, ZN => gl_rom_n_1222);
  gl_rom_g35199 : ND4D0BWP7T port map(A1 => gl_rom_n_660, A2 => gl_rom_n_664, A3 => gl_rom_n_668, A4 => gl_rom_n_657, ZN => gl_rom_n_1221);
  gl_rom_g35200 : ND4D0BWP7T port map(A1 => gl_rom_n_665, A2 => gl_rom_n_655, A3 => gl_rom_n_663, A4 => gl_rom_n_648, ZN => gl_rom_n_1220);
  gl_rom_g35201 : ND4D0BWP7T port map(A1 => gl_rom_n_659, A2 => gl_rom_n_661, A3 => gl_rom_n_662, A4 => gl_rom_n_658, ZN => gl_rom_n_1219);
  gl_rom_g35202 : ND4D0BWP7T port map(A1 => gl_rom_n_645, A2 => gl_rom_n_650, A3 => gl_rom_n_653, A4 => gl_rom_n_643, ZN => gl_rom_n_1218);
  gl_rom_g35203 : ND4D0BWP7T port map(A1 => gl_rom_n_654, A2 => gl_rom_n_656, A3 => gl_rom_n_651, A4 => gl_rom_n_649, ZN => gl_rom_n_1217);
  gl_rom_g35204 : ND4D0BWP7T port map(A1 => gl_rom_n_647, A2 => gl_rom_n_644, A3 => gl_rom_n_646, A4 => gl_rom_n_642, ZN => gl_rom_n_1216);
  gl_rom_g35205 : ND4D0BWP7T port map(A1 => gl_rom_n_638, A2 => gl_rom_n_640, A3 => gl_rom_n_635, A4 => gl_rom_n_634, ZN => gl_rom_n_1215);
  gl_rom_g35206 : ND4D0BWP7T port map(A1 => gl_rom_n_589, A2 => gl_rom_n_628, A3 => gl_rom_n_623, A4 => gl_rom_n_608, ZN => gl_rom_n_1214);
  gl_rom_g35207 : ND4D0BWP7T port map(A1 => gl_rom_n_627, A2 => gl_rom_n_637, A3 => gl_rom_n_633, A4 => gl_rom_n_630, ZN => gl_rom_n_1213);
  gl_rom_g35208 : ND4D0BWP7T port map(A1 => gl_rom_n_619, A2 => gl_rom_n_632, A3 => gl_rom_n_624, A4 => gl_rom_n_616, ZN => gl_rom_n_1212);
  gl_rom_g35209 : ND4D0BWP7T port map(A1 => gl_rom_n_625, A2 => gl_rom_n_631, A3 => gl_rom_n_629, A4 => gl_rom_n_626, ZN => gl_rom_n_1211);
  gl_rom_g35210 : ND4D0BWP7T port map(A1 => gl_rom_n_617, A2 => gl_rom_n_620, A3 => gl_rom_n_622, A4 => gl_rom_n_615, ZN => gl_rom_n_1210);
  gl_rom_g35211 : ND4D0BWP7T port map(A1 => gl_rom_n_609, A2 => gl_rom_n_621, A3 => gl_rom_n_618, A4 => gl_rom_n_614, ZN => gl_rom_n_1209);
  gl_rom_g35212 : ND4D0BWP7T port map(A1 => gl_rom_n_611, A2 => gl_rom_n_612, A3 => gl_rom_n_613, A4 => gl_rom_n_610, ZN => gl_rom_n_1208);
  gl_rom_g35213 : ND4D0BWP7T port map(A1 => gl_rom_n_596, A2 => gl_rom_n_581, A3 => gl_rom_n_600, A4 => gl_rom_n_588, ZN => gl_rom_n_1207);
  gl_rom_g35214 : ND4D0BWP7T port map(A1 => gl_rom_n_603, A2 => gl_rom_n_606, A3 => gl_rom_n_607, A4 => gl_rom_n_602, ZN => gl_rom_n_1206);
  gl_rom_g35215 : ND4D0BWP7T port map(A1 => gl_rom_n_605, A2 => gl_rom_n_598, A3 => gl_rom_n_601, A4 => gl_rom_n_593, ZN => gl_rom_n_1205);
  gl_rom_g35216 : ND4D0BWP7T port map(A1 => gl_rom_n_597, A2 => gl_rom_n_599, A3 => gl_rom_n_595, A4 => gl_rom_n_594, ZN => gl_rom_n_1204);
  gl_rom_g35217 : ND4D0BWP7T port map(A1 => gl_rom_n_585, A2 => gl_rom_n_579, A3 => gl_rom_n_591, A4 => gl_rom_n_584, ZN => gl_rom_n_1203);
  gl_rom_g35218 : ND4D0BWP7T port map(A1 => gl_rom_n_590, A2 => gl_rom_n_592, A3 => gl_rom_n_587, A4 => gl_rom_n_586, ZN => gl_rom_n_1202);
  gl_rom_g35219 : ND4D0BWP7T port map(A1 => gl_rom_n_582, A2 => gl_rom_n_583, A3 => gl_rom_n_580, A4 => gl_rom_n_578, ZN => gl_rom_n_1201);
  gl_rom_g35220 : ND4D0BWP7T port map(A1 => gl_rom_n_455, A2 => gl_rom_n_604, A3 => gl_rom_n_577, A4 => gl_rom_n_482, ZN => gl_rom_n_1200);
  gl_rom_g35221 : ND4D0BWP7T port map(A1 => gl_rom_n_514, A2 => gl_rom_n_575, A3 => gl_rom_n_545, A4 => gl_rom_n_490, ZN => gl_rom_n_1199);
  gl_rom_g35222 : ND4D0BWP7T port map(A1 => gl_rom_n_572, A2 => gl_rom_n_573, A3 => gl_rom_n_576, A4 => gl_rom_n_569, ZN => gl_rom_n_1198);
  gl_rom_g35223 : ND4D0BWP7T port map(A1 => gl_rom_n_568, A2 => gl_rom_n_542, A3 => gl_rom_n_558, A4 => gl_rom_n_529, ZN => gl_rom_n_1197);
  gl_rom_g35224 : ND4D0BWP7T port map(A1 => gl_rom_n_574, A2 => gl_rom_n_566, A3 => gl_rom_n_570, A4 => gl_rom_n_564, ZN => gl_rom_n_1196);
  gl_rom_g35225 : ND4D0BWP7T port map(A1 => gl_rom_n_554, A2 => gl_rom_n_561, A3 => gl_rom_n_571, A4 => gl_rom_n_551, ZN => gl_rom_n_1195);
  gl_rom_g35226 : ND4D0BWP7T port map(A1 => gl_rom_n_565, A2 => gl_rom_n_567, A3 => gl_rom_n_563, A4 => gl_rom_n_562, ZN => gl_rom_n_1194);
  gl_rom_g35227 : ND4D0BWP7T port map(A1 => gl_rom_n_556, A2 => gl_rom_n_548, A3 => gl_rom_n_560, A4 => gl_rom_n_552, ZN => gl_rom_n_1193);
  gl_rom_g35228 : ND4D0BWP7T port map(A1 => gl_rom_n_557, A2 => gl_rom_n_559, A3 => gl_rom_n_555, A4 => gl_rom_n_553, ZN => gl_rom_n_1192);
  gl_rom_g35229 : ND4D0BWP7T port map(A1 => gl_rom_n_911, A2 => gl_rom_n_756, A3 => gl_rom_n_862, A4 => gl_rom_n_641, ZN => gl_rom_n_1191);
  gl_rom_g35230 : ND4D0BWP7T port map(A1 => gl_rom_n_39, A2 => gl_rom_n_41, A3 => gl_rom_n_43, A4 => gl_rom_n_806, ZN => gl_rom_n_1190);
  gl_rom_g35231 : ND4D0BWP7T port map(A1 => gl_rom_n_543, A2 => gl_rom_n_544, A3 => gl_rom_n_539, A4 => gl_rom_n_537, ZN => gl_rom_n_1189);
  gl_rom_g35232 : ND4D0BWP7T port map(A1 => gl_rom_n_535, A2 => gl_rom_n_538, A3 => gl_rom_n_541, A4 => gl_rom_n_531, ZN => gl_rom_n_1188);
  gl_rom_g35233 : ND4D0BWP7T port map(A1 => gl_rom_n_534, A2 => gl_rom_n_530, A3 => gl_rom_n_536, A4 => gl_rom_n_532, ZN => gl_rom_n_1187);
  gl_rom_g35234 : ND4D0BWP7T port map(A1 => gl_rom_n_528, A2 => gl_rom_n_523, A3 => gl_rom_n_526, A4 => gl_rom_n_522, ZN => gl_rom_n_1186);
  gl_rom_g35235 : ND4D0BWP7T port map(A1 => gl_rom_n_517, A2 => gl_rom_n_525, A3 => gl_rom_n_524, A4 => gl_rom_n_519, ZN => gl_rom_n_1185);
  gl_rom_g35236 : ND4D0BWP7T port map(A1 => gl_rom_n_521, A2 => gl_rom_n_516, A3 => gl_rom_n_518, A4 => gl_rom_n_515, ZN => gl_rom_n_1184);
  gl_rom_g35237 : ND4D0BWP7T port map(A1 => gl_rom_n_498, A2 => gl_rom_n_476, A3 => gl_rom_n_510, A4 => gl_rom_n_480, ZN => gl_rom_n_1183);
  gl_rom_g35238 : ND4D0BWP7T port map(A1 => gl_rom_n_509, A2 => gl_rom_n_512, A3 => gl_rom_n_513, A4 => gl_rom_n_508, ZN => gl_rom_n_1182);
  gl_rom_g35239 : ND4D0BWP7T port map(A1 => gl_rom_n_511, A2 => gl_rom_n_504, A3 => gl_rom_n_507, A4 => gl_rom_n_501, ZN => gl_rom_n_1181);
  gl_rom_g35240 : ND4D0BWP7T port map(A1 => gl_rom_n_487, A2 => gl_rom_n_505, A3 => gl_rom_n_502, A4 => gl_rom_n_493, ZN => gl_rom_n_1180);
  gl_rom_g35241 : ND4D0BWP7T port map(A1 => gl_rom_n_500, A2 => gl_rom_n_503, A3 => gl_rom_n_506, A4 => gl_rom_n_499, ZN => gl_rom_n_1179);
  gl_rom_g35242 : ND4D0BWP7T port map(A1 => gl_rom_n_425, A2 => gl_rom_n_271, A3 => gl_rom_n_326, A4 => gl_rom_n_203, ZN => gl_rom_n_1178);
  gl_rom_g35243 : ND4D0BWP7T port map(A1 => gl_rom_n_488, A2 => gl_rom_n_492, A3 => gl_rom_n_496, A4 => gl_rom_n_485, ZN => gl_rom_n_1177);
  gl_rom_g35244 : ND4D0BWP7T port map(A1 => gl_rom_n_495, A2 => gl_rom_n_497, A3 => gl_rom_n_494, A4 => gl_rom_n_491, ZN => gl_rom_n_1176);
  gl_rom_g35245 : ND4D0BWP7T port map(A1 => gl_rom_n_484, A2 => gl_rom_n_486, A3 => gl_rom_n_489, A4 => gl_rom_n_483, ZN => gl_rom_n_1175);
  gl_rom_g35246 : ND4D0BWP7T port map(A1 => gl_rom_n_477, A2 => gl_rom_n_479, A3 => gl_rom_n_481, A4 => gl_rom_n_474, ZN => gl_rom_n_1174);
  gl_rom_g35247 : ND4D0BWP7T port map(A1 => gl_rom_n_478, A2 => gl_rom_n_469, A3 => gl_rom_n_475, A4 => gl_rom_n_467, ZN => gl_rom_n_1173);
  gl_rom_g35248 : ND4D0BWP7T port map(A1 => gl_rom_n_462, A2 => gl_rom_n_473, A3 => gl_rom_n_471, A4 => gl_rom_n_454, ZN => gl_rom_n_1172);
  gl_rom_g35249 : ND4D0BWP7T port map(A1 => gl_rom_n_466, A2 => gl_rom_n_472, A3 => gl_rom_n_470, A4 => gl_rom_n_468, ZN => gl_rom_n_1171);
  gl_rom_g35250 : ND4D0BWP7T port map(A1 => gl_rom_n_419, A2 => gl_rom_n_363, A3 => gl_rom_n_450, A4 => gl_rom_n_386, ZN => gl_rom_n_1170);
  gl_rom_g35251 : ND4D0BWP7T port map(A1 => gl_rom_n_464, A2 => gl_rom_n_457, A3 => gl_rom_n_460, A4 => gl_rom_n_452, ZN => gl_rom_n_1169);
  gl_rom_g35252 : ND4D0BWP7T port map(A1 => gl_rom_n_463, A2 => gl_rom_n_459, A3 => gl_rom_n_465, A4 => gl_rom_n_461, ZN => gl_rom_n_1168);
  gl_rom_g35253 : ND4D0BWP7T port map(A1 => gl_rom_n_458, A2 => gl_rom_n_453, A3 => gl_rom_n_456, A4 => gl_rom_n_451, ZN => gl_rom_n_1167);
  gl_rom_g35254 : ND4D0BWP7T port map(A1 => gl_rom_n_443, A2 => gl_rom_n_449, A3 => gl_rom_n_447, A4 => gl_rom_n_446, ZN => gl_rom_n_1166);
  gl_rom_g35255 : ND4D0BWP7T port map(A1 => gl_rom_n_401, A2 => gl_rom_n_445, A3 => gl_rom_n_432, A4 => gl_rom_n_416, ZN => gl_rom_n_1165);
  gl_rom_g35256 : ND4D0BWP7T port map(A1 => gl_rom_n_448, A2 => gl_rom_n_440, A3 => gl_rom_n_444, A4 => gl_rom_n_438, ZN => gl_rom_n_1164);
  gl_rom_g35257 : ND4D0BWP7T port map(A1 => gl_rom_n_435, A2 => gl_rom_n_424, A3 => gl_rom_n_442, A4 => gl_rom_n_428, ZN => gl_rom_n_1163);
  gl_rom_g35258 : ND4D0BWP7T port map(A1 => gl_rom_n_437, A2 => gl_rom_n_439, A3 => gl_rom_n_441, A4 => gl_rom_n_436, ZN => gl_rom_n_1162);
  gl_rom_g35259 : ND4D0BWP7T port map(A1 => gl_rom_n_430, A2 => gl_rom_n_434, A3 => gl_rom_n_426, A4 => gl_rom_n_421, ZN => gl_rom_n_1161);
  gl_rom_g35260 : ND4D0BWP7T port map(A1 => gl_rom_n_429, A2 => gl_rom_n_431, A3 => gl_rom_n_433, A4 => gl_rom_n_427, ZN => gl_rom_n_1160);
  gl_rom_g35261 : ND4D0BWP7T port map(A1 => gl_rom_n_420, A2 => gl_rom_n_422, A3 => gl_rom_n_423, A4 => gl_rom_n_418, ZN => gl_rom_n_1159);
  gl_rom_g35262 : ND4D0BWP7T port map(A1 => gl_rom_n_413, A2 => gl_rom_n_415, A3 => gl_rom_n_417, A4 => gl_rom_n_411, ZN => gl_rom_n_1158);
  gl_rom_g35263 : ND4D0BWP7T port map(A1 => gl_rom_n_410, A2 => gl_rom_n_414, A3 => gl_rom_n_407, A4 => gl_rom_n_406, ZN => gl_rom_n_1157);
  gl_rom_g35264 : ND4D0BWP7T port map(A1 => gl_rom_n_398, A2 => gl_rom_n_412, A3 => gl_rom_n_403, A4 => gl_rom_n_393, ZN => gl_rom_n_1156);
  gl_rom_g35265 : ND4D0BWP7T port map(A1 => gl_rom_n_409, A2 => gl_rom_n_405, A3 => gl_rom_n_408, A4 => gl_rom_n_404, ZN => gl_rom_n_1155);
  gl_rom_g35266 : ND4D0BWP7T port map(A1 => gl_rom_n_397, A2 => gl_rom_n_399, A3 => gl_rom_n_402, A4 => gl_rom_n_395, ZN => gl_rom_n_1154);
  gl_rom_g35267 : ND4D0BWP7T port map(A1 => gl_rom_n_392, A2 => gl_rom_n_396, A3 => gl_rom_n_400, A4 => gl_rom_n_390, ZN => gl_rom_n_1153);
  gl_rom_g35268 : ND4D0BWP7T port map(A1 => gl_rom_n_394, A2 => gl_rom_n_389, A3 => gl_rom_n_391, A4 => gl_rom_n_388, ZN => gl_rom_n_1152);
  gl_rom_g35269 : ND4D0BWP7T port map(A1 => gl_rom_n_370, A2 => gl_rom_n_384, A3 => gl_rom_n_353, A4 => gl_rom_n_342, ZN => gl_rom_n_1151);
  gl_rom_g35270 : ND4D0BWP7T port map(A1 => gl_rom_n_381, A2 => gl_rom_n_383, A3 => gl_rom_n_385, A4 => gl_rom_n_379, ZN => gl_rom_n_1150);
  gl_rom_g35271 : ND4D0BWP7T port map(A1 => gl_rom_n_382, A2 => gl_rom_n_376, A3 => gl_rom_n_380, A4 => gl_rom_n_373, ZN => gl_rom_n_1149);
  gl_rom_g35272 : ND4D0BWP7T port map(A1 => gl_rom_n_378, A2 => gl_rom_n_362, A3 => gl_rom_n_374, A4 => gl_rom_n_359, ZN => gl_rom_n_1148);
  gl_rom_g35273 : ND4D0BWP7T port map(A1 => gl_rom_n_372, A2 => gl_rom_n_375, A3 => gl_rom_n_377, A4 => gl_rom_n_371, ZN => gl_rom_n_1147);
  gl_rom_g35274 : ND4D0BWP7T port map(A1 => gl_rom_n_357, A2 => gl_rom_n_368, A3 => gl_rom_n_365, A4 => gl_rom_n_361, ZN => gl_rom_n_1146);
  gl_rom_g35275 : ND4D0BWP7T port map(A1 => gl_rom_n_366, A2 => gl_rom_n_367, A3 => gl_rom_n_369, A4 => gl_rom_n_364, ZN => gl_rom_n_1145);
  gl_rom_g35276 : ND4D0BWP7T port map(A1 => gl_rom_n_356, A2 => gl_rom_n_358, A3 => gl_rom_n_360, A4 => gl_rom_n_355, ZN => gl_rom_n_1144);
  gl_rom_g35277 : ND4D0BWP7T port map(A1 => gl_rom_n_329, A2 => gl_rom_n_350, A3 => gl_rom_n_341, A4 => gl_rom_n_331, ZN => gl_rom_n_1143);
  gl_rom_g35278 : ND4D0BWP7T port map(A1 => gl_rom_n_349, A2 => gl_rom_n_351, A3 => gl_rom_n_354, A4 => gl_rom_n_347, ZN => gl_rom_n_1142);
  gl_rom_g35279 : ND4D0BWP7T port map(A1 => gl_rom_n_348, A2 => gl_rom_n_339, A3 => gl_rom_n_352, A4 => gl_rom_n_343, ZN => gl_rom_n_1141);
  gl_rom_g35280 : ND4D0BWP7T port map(A1 => gl_rom_n_338, A2 => gl_rom_n_346, A3 => gl_rom_n_344, A4 => gl_rom_n_340, ZN => gl_rom_n_1140);
  gl_rom_g35281 : ND4D0BWP7T port map(A1 => gl_rom_n_257, A2 => gl_rom_n_345, A3 => gl_rom_n_289, A4 => gl_rom_n_265, ZN => gl_rom_n_1139);
  gl_rom_g35282 : ND4D0BWP7T port map(A1 => gl_rom_n_336, A2 => gl_rom_n_328, A3 => gl_rom_n_334, A4 => gl_rom_n_325, ZN => gl_rom_n_1138);
  gl_rom_g35283 : ND4D0BWP7T port map(A1 => gl_rom_n_333, A2 => gl_rom_n_335, A3 => gl_rom_n_337, A4 => gl_rom_n_332, ZN => gl_rom_n_1137);
  gl_rom_g35284 : ND4D0BWP7T port map(A1 => gl_rom_n_327, A2 => gl_rom_n_330, A3 => gl_rom_n_324, A4 => gl_rom_n_323, ZN => gl_rom_n_1136);
  gl_rom_g35285 : ND4D0BWP7T port map(A1 => gl_rom_n_288, A2 => gl_rom_n_302, A3 => gl_rom_n_322, A4 => gl_rom_n_279, ZN => gl_rom_n_1135);
  gl_rom_g35286 : ND4D0BWP7T port map(A1 => gl_rom_n_315, A2 => gl_rom_n_321, A3 => gl_rom_n_319, A4 => gl_rom_n_318, ZN => gl_rom_n_1134);
  gl_rom_g35287 : ND4D0BWP7T port map(A1 => gl_rom_n_317, A2 => gl_rom_n_298, A3 => gl_rom_n_309, A4 => gl_rom_n_293, ZN => gl_rom_n_1133);
  gl_rom_g35288 : ND4D0BWP7T port map(A1 => gl_rom_n_312, A2 => gl_rom_n_316, A3 => gl_rom_n_320, A4 => gl_rom_n_308, ZN => gl_rom_n_1132);
  gl_rom_g35289 : ND4D0BWP7T port map(A1 => gl_rom_n_304, A2 => gl_rom_n_313, A3 => gl_rom_n_314, A4 => gl_rom_n_301, ZN => gl_rom_n_1131);
  gl_rom_g35290 : ND4D0BWP7T port map(A1 => gl_rom_n_310, A2 => gl_rom_n_311, A3 => gl_rom_n_307, A4 => gl_rom_n_306, ZN => gl_rom_n_1130);
  gl_rom_g35291 : ND4D0BWP7T port map(A1 => gl_rom_n_299, A2 => gl_rom_n_305, A3 => gl_rom_n_303, A4 => gl_rom_n_300, ZN => gl_rom_n_1129);
  gl_rom_g35292 : ND4D0BWP7T port map(A1 => gl_rom_n_286, A2 => gl_rom_n_297, A3 => gl_rom_n_296, A4 => gl_rom_n_291, ZN => gl_rom_n_1128);
  gl_rom_g35293 : ND4D0BWP7T port map(A1 => gl_rom_n_292, A2 => gl_rom_n_550, A3 => gl_rom_n_295, A4 => gl_rom_n_290, ZN => gl_rom_n_1127);
  gl_rom_g35294 : ND4D0BWP7T port map(A1 => gl_rom_n_284, A2 => gl_rom_n_285, A3 => gl_rom_n_287, A4 => gl_rom_n_283, ZN => gl_rom_n_1126);
  gl_rom_g35295 : ND4D0BWP7T port map(A1 => gl_rom_n_282, A2 => gl_rom_n_270, A3 => gl_rom_n_281, A4 => gl_rom_n_262, ZN => gl_rom_n_1125);
  gl_rom_g35296 : ND4D0BWP7T port map(A1 => gl_rom_n_276, A2 => gl_rom_n_278, A3 => gl_rom_n_280, A4 => gl_rom_n_274, ZN => gl_rom_n_1124);
  gl_rom_g35297 : ND4D0BWP7T port map(A1 => gl_rom_n_275, A2 => gl_rom_n_277, A3 => gl_rom_n_269, A4 => gl_rom_n_266, ZN => gl_rom_n_1123);
  gl_rom_g35298 : ND4D0BWP7T port map(A1 => gl_rom_n_268, A2 => gl_rom_n_272, A3 => gl_rom_n_273, A4 => gl_rom_n_267, ZN => gl_rom_n_1122);
  gl_rom_g35299 : ND4D0BWP7T port map(A1 => gl_rom_n_254, A2 => gl_rom_n_259, A3 => gl_rom_n_261, A4 => gl_rom_n_250, ZN => gl_rom_n_1121);
  gl_rom_g35300 : ND4D0BWP7T port map(A1 => gl_rom_n_260, A2 => gl_rom_n_263, A3 => gl_rom_n_264, A4 => gl_rom_n_258, ZN => gl_rom_n_1120);
  gl_rom_g35301 : ND4D0BWP7T port map(A1 => gl_rom_n_252, A2 => gl_rom_n_255, A3 => gl_rom_n_256, A4 => gl_rom_n_251, ZN => gl_rom_n_1119);
  gl_rom_g35302 : ND4D0BWP7T port map(A1 => gl_rom_n_218, A2 => gl_rom_n_253, A3 => gl_rom_n_249, A4 => gl_rom_n_223, ZN => gl_rom_n_1118);
  gl_rom_g35303 : ND4D0BWP7T port map(A1 => gl_rom_n_243, A2 => gl_rom_n_248, A3 => gl_rom_n_247, A4 => gl_rom_n_245, ZN => gl_rom_n_1117);
  gl_rom_g35304 : ND4D0BWP7T port map(A1 => gl_rom_n_239, A2 => gl_rom_n_242, A3 => gl_rom_n_246, A4 => gl_rom_n_237, ZN => gl_rom_n_1116);
  gl_rom_g35305 : ND4D0BWP7T port map(A1 => gl_rom_n_235, A2 => gl_rom_n_227, A3 => gl_rom_n_244, A4 => gl_rom_n_231, ZN => gl_rom_n_1115);
  gl_rom_g35306 : ND4D0BWP7T port map(A1 => gl_rom_n_236, A2 => gl_rom_n_241, A3 => gl_rom_n_240, A4 => gl_rom_n_238, ZN => gl_rom_n_1114);
  gl_rom_g35307 : ND4D0BWP7T port map(A1 => gl_rom_n_228, A2 => gl_rom_n_232, A3 => gl_rom_n_225, A4 => gl_rom_n_222, ZN => gl_rom_n_1113);
  gl_rom_g35308 : ND4D0BWP7T port map(A1 => gl_rom_n_229, A2 => gl_rom_n_234, A3 => gl_rom_n_233, A4 => gl_rom_n_230, ZN => gl_rom_n_1112);
  gl_rom_g35309 : ND4D0BWP7T port map(A1 => gl_rom_n_220, A2 => gl_rom_n_226, A3 => gl_rom_n_224, A4 => gl_rom_n_221, ZN => gl_rom_n_1111);
  gl_rom_g35310 : ND4D0BWP7T port map(A1 => gl_rom_n_217, A2 => gl_rom_n_219, A3 => gl_rom_n_214, A4 => gl_rom_n_213, ZN => gl_rom_n_1110);
  gl_rom_g35311 : ND4D0BWP7T port map(A1 => gl_rom_n_216, A2 => gl_rom_n_199, A3 => gl_rom_n_211, A4 => gl_rom_n_193, ZN => gl_rom_n_1109);
  gl_rom_g35312 : ND4D0BWP7T port map(A1 => gl_rom_n_195, A2 => gl_rom_n_144, A3 => gl_rom_n_180, A4 => gl_rom_n_116, ZN => gl_rom_n_1108);
  gl_rom_g35313 : ND4D0BWP7T port map(A1 => gl_rom_n_208, A2 => gl_rom_n_212, A3 => gl_rom_n_215, A4 => gl_rom_n_205, ZN => gl_rom_n_1107);
  gl_rom_g35314 : ND4D0BWP7T port map(A1 => gl_rom_n_207, A2 => gl_rom_n_210, A3 => gl_rom_n_209, A4 => gl_rom_n_206, ZN => gl_rom_n_1106);
  gl_rom_g35315 : ND4D0BWP7T port map(A1 => gl_rom_n_189, A2 => gl_rom_n_201, A3 => gl_rom_n_197, A4 => gl_rom_n_191, ZN => gl_rom_n_1105);
  gl_rom_g35316 : ND4D0BWP7T port map(A1 => gl_rom_n_204, A2 => gl_rom_n_198, A3 => gl_rom_n_200, A4 => gl_rom_n_196, ZN => gl_rom_n_1104);
  gl_rom_g35317 : ND4D0BWP7T port map(A1 => gl_rom_n_192, A2 => gl_rom_n_188, A3 => gl_rom_n_194, A4 => gl_rom_n_190, ZN => gl_rom_n_1103);
  gl_rom_g35318 : ND4D0BWP7T port map(A1 => gl_rom_n_184, A2 => gl_rom_n_186, A3 => gl_rom_n_187, A4 => gl_rom_n_181, ZN => gl_rom_n_1102);
  gl_rom_g35319 : ND4D0BWP7T port map(A1 => gl_rom_n_178, A2 => gl_rom_n_163, A3 => gl_rom_n_183, A4 => gl_rom_n_169, ZN => gl_rom_n_1101);
  gl_rom_g35320 : ND4D0BWP7T port map(A1 => gl_rom_n_176, A2 => gl_rom_n_182, A3 => gl_rom_n_185, A4 => gl_rom_n_172, ZN => gl_rom_n_1100);
  gl_rom_g35321 : ND4D0BWP7T port map(A1 => gl_rom_n_140, A2 => gl_rom_n_175, A3 => gl_rom_n_171, A4 => gl_rom_n_151, ZN => gl_rom_n_1099);
  gl_rom_g35322 : ND4D0BWP7T port map(A1 => gl_rom_n_173, A2 => gl_rom_n_179, A3 => gl_rom_n_177, A4 => gl_rom_n_174, ZN => gl_rom_n_1098);
  gl_rom_g35323 : ND4D0BWP7T port map(A1 => gl_rom_n_165, A2 => gl_rom_n_170, A3 => gl_rom_n_167, A4 => gl_rom_n_164, ZN => gl_rom_n_1097);
  gl_rom_g35324 : ND4D0BWP7T port map(A1 => gl_rom_n_162, A2 => gl_rom_n_166, A3 => gl_rom_n_168, A4 => gl_rom_n_159, ZN => gl_rom_n_1096);
  gl_rom_g35325 : ND4D0BWP7T port map(A1 => gl_rom_n_161, A2 => gl_rom_n_158, A3 => gl_rom_n_160, A4 => gl_rom_n_157, ZN => gl_rom_n_1095);
  gl_rom_g35326 : ND4D0BWP7T port map(A1 => gl_rom_n_154, A2 => gl_rom_n_139, A3 => gl_rom_n_148, A4 => gl_rom_n_132, ZN => gl_rom_n_1094);
  gl_rom_g35327 : ND4D0BWP7T port map(A1 => gl_rom_n_152, A2 => gl_rom_n_156, A3 => gl_rom_n_155, A4 => gl_rom_n_150, ZN => gl_rom_n_1093);
  gl_rom_g35328 : ND4D0BWP7T port map(A1 => gl_rom_n_145, A2 => gl_rom_n_149, A3 => gl_rom_n_153, A4 => gl_rom_n_141, ZN => gl_rom_n_1092);
  gl_rom_g35329 : ND4D0BWP7T port map(A1 => gl_rom_n_142, A2 => gl_rom_n_147, A3 => gl_rom_n_146, A4 => gl_rom_n_143, ZN => gl_rom_n_1091);
  gl_rom_g35330 : ND4D0BWP7T port map(A1 => gl_rom_n_127, A2 => gl_rom_n_136, A3 => gl_rom_n_134, A4 => gl_rom_n_130, ZN => gl_rom_n_1090);
  gl_rom_g35331 : ND4D0BWP7T port map(A1 => gl_rom_n_138, A2 => gl_rom_n_135, A3 => gl_rom_n_137, A4 => gl_rom_n_133, ZN => gl_rom_n_1089);
  gl_rom_g35332 : ND4D0BWP7T port map(A1 => gl_rom_n_131, A2 => gl_rom_n_128, A3 => gl_rom_n_129, A4 => gl_rom_n_126, ZN => gl_rom_n_1088);
  gl_rom_g35333 : ND4D0BWP7T port map(A1 => gl_rom_n_93, A2 => gl_rom_n_1028, A3 => gl_rom_n_72, A4 => gl_rom_n_973, ZN => gl_rom_n_1087);
  gl_rom_g35334 : ND4D0BWP7T port map(A1 => gl_rom_n_125, A2 => gl_rom_n_121, A3 => gl_rom_n_124, A4 => gl_rom_n_120, ZN => gl_rom_n_1086);
  gl_rom_g35335 : ND4D0BWP7T port map(A1 => gl_rom_n_78, A2 => gl_rom_n_387, A3 => gl_rom_n_772, A4 => gl_rom_n_202, ZN => gl_rom_n_1085);
  gl_rom_g35336 : ND4D0BWP7T port map(A1 => gl_rom_n_75, A2 => gl_rom_n_119, A3 => gl_rom_n_109, A4 => gl_rom_n_91, ZN => gl_rom_n_1084);
  gl_rom_g35337 : ND4D0BWP7T port map(A1 => gl_rom_n_101, A2 => gl_rom_n_122, A3 => gl_rom_n_114, A4 => gl_rom_n_107, ZN => gl_rom_n_1083);
  gl_rom_g35338 : ND4D0BWP7T port map(A1 => gl_rom_n_113, A2 => gl_rom_n_118, A3 => gl_rom_n_123, A4 => gl_rom_n_112, ZN => gl_rom_n_1082);
  gl_rom_g35339 : ND4D0BWP7T port map(A1 => gl_rom_n_115, A2 => gl_rom_n_110, A3 => gl_rom_n_117, A4 => gl_rom_n_111, ZN => gl_rom_n_1081);
  gl_rom_g35340 : ND4D0BWP7T port map(A1 => gl_rom_n_99, A2 => gl_rom_n_104, A3 => gl_rom_n_106, A4 => gl_rom_n_97, ZN => gl_rom_n_1080);
  gl_rom_g35341 : ND4D0BWP7T port map(A1 => gl_rom_n_105, A2 => gl_rom_n_108, A3 => gl_rom_n_103, A4 => gl_rom_n_102, ZN => gl_rom_n_1079);
  gl_rom_g35342 : ND4D0BWP7T port map(A1 => gl_rom_n_96, A2 => gl_rom_n_100, A3 => gl_rom_n_98, A4 => gl_rom_n_95, ZN => gl_rom_n_1078);
  gl_rom_g35343 : ND4D0BWP7T port map(A1 => gl_rom_n_88, A2 => gl_rom_n_92, A3 => gl_rom_n_94, A4 => gl_rom_n_87, ZN => gl_rom_n_1077);
  gl_rom_g35344 : ND4D0BWP7T port map(A1 => gl_rom_n_89, A2 => gl_rom_n_77, A3 => gl_rom_n_85, A4 => gl_rom_n_68, ZN => gl_rom_n_1076);
  gl_rom_g35345 : ND4D0BWP7T port map(A1 => gl_rom_n_82, A2 => gl_rom_n_86, A3 => gl_rom_n_90, A4 => gl_rom_n_79, ZN => gl_rom_n_1075);
  gl_rom_g35346 : ND4D0BWP7T port map(A1 => gl_rom_n_81, A2 => gl_rom_n_83, A3 => gl_rom_n_84, A4 => gl_rom_n_80, ZN => gl_rom_n_1074);
  gl_rom_g35347 : ND4D0BWP7T port map(A1 => gl_rom_n_65, A2 => gl_rom_n_70, A3 => gl_rom_n_74, A4 => gl_rom_n_63, ZN => gl_rom_n_1073);
  gl_rom_g35348 : ND4D0BWP7T port map(A1 => gl_rom_n_73, A2 => gl_rom_n_76, A3 => gl_rom_n_71, A4 => gl_rom_n_69, ZN => gl_rom_n_1072);
  gl_rom_g35349 : ND4D0BWP7T port map(A1 => gl_rom_n_64, A2 => gl_rom_n_66, A3 => gl_rom_n_67, A4 => gl_rom_n_62, ZN => gl_rom_n_1071);
  gl_rom_g35350 : ND4D0BWP7T port map(A1 => gl_rom_n_55, A2 => gl_rom_n_61, A3 => gl_rom_n_60, A4 => gl_rom_n_57, ZN => gl_rom_n_1070);
  gl_rom_g35351 : ND4D0BWP7T port map(A1 => gl_rom_n_58, A2 => gl_rom_n_44, A3 => gl_rom_n_53, A4 => gl_rom_n_1055, ZN => gl_rom_n_1069);
  gl_rom_g35352 : ND4D0BWP7T port map(A1 => gl_rom_n_52, A2 => gl_rom_n_56, A3 => gl_rom_n_59, A4 => gl_rom_n_49, ZN => gl_rom_n_1068);
  gl_rom_g35353 : ND4D0BWP7T port map(A1 => gl_rom_n_1053, A2 => gl_rom_n_50, A3 => gl_rom_n_45, A4 => gl_rom_n_1042, ZN => gl_rom_n_1067);
  gl_rom_g35354 : ND4D0BWP7T port map(A1 => gl_rom_n_48, A2 => gl_rom_n_51, A3 => gl_rom_n_54, A4 => gl_rom_n_47, ZN => gl_rom_n_1066);
  gl_rom_g35355 : ND4D0BWP7T port map(A1 => gl_rom_n_46, A2 => gl_rom_n_1021, A3 => gl_rom_n_1054, A4 => gl_rom_n_988, ZN => gl_rom_n_1065);
  gl_rom_g35356 : ND4D0BWP7T port map(A1 => gl_rom_n_1061, A2 => gl_rom_n_40, A3 => gl_rom_n_42, A4 => gl_rom_n_1058, ZN => gl_rom_n_1064);
  gl_rom_g35357 : ND4D0BWP7T port map(A1 => gl_rom_n_527, A2 => gl_rom_n_540, A3 => gl_rom_n_533, A4 => gl_rom_n_520, ZN => gl_rom_n_1063);
  gl_rom_g35358 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_776(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_779(0), ZN => gl_rom_n_1062);
  gl_rom_g35359 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_385(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_389(0), ZN => gl_rom_n_1061);
  gl_rom_g35360 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_977(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_981(1), ZN => gl_rom_n_1060);
  gl_rom_g35361 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_980(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_982(1), ZN => gl_rom_n_1059);
  gl_rom_g35362 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_384(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_387(0), ZN => gl_rom_n_1058);
  gl_rom_g35363 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_978(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_979(1), ZN => gl_rom_n_1057);
  gl_rom_g35364 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_976(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_983(1), ZN => gl_rom_n_1056);
  gl_rom_g35365 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_712(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_713(0), ZN => gl_rom_n_1055);
  gl_rom_g35366 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_956(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_958(0), ZN => gl_rom_n_1054);
  gl_rom_g35367 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_882(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_887(0), ZN => gl_rom_n_1053);
  gl_rom_g35368 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_706(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_711(0), ZN => gl_rom_n_1052);
  gl_rom_g35369 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_985(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_989(1), ZN => gl_rom_n_1051);
  gl_rom_g35370 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_988(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_990(1), ZN => gl_rom_n_1050);
  gl_rom_g35371 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_378(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_383(0), ZN => gl_rom_n_1049);
  gl_rom_g35372 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_986(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_987(1), ZN => gl_rom_n_1048);
  gl_rom_g35373 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_984(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_991(1), ZN => gl_rom_n_1047);
  gl_rom_g35374 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_708(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_710(0), ZN => gl_rom_n_1046);
  gl_rom_g35375 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_380(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_382(0), ZN => gl_rom_n_1045);
  gl_rom_g35376 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_994(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_999(1), ZN => gl_rom_n_1044);
  gl_rom_g35377 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_993(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_997(1), ZN => gl_rom_n_1043);
  gl_rom_g35378 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_880(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_883(0), ZN => gl_rom_n_1042);
  gl_rom_g35379 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_381(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_379(0), ZN => gl_rom_n_1041);
  gl_rom_g35380 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_996(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_998(1), ZN => gl_rom_n_1040);
  gl_rom_g35381 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_376(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_377(0), ZN => gl_rom_n_1039);
  gl_rom_g35382 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_992(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_995(1), ZN => gl_rom_n_1038);
  gl_rom_g35383 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_1022(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_1023(1), ZN => gl_rom_n_1037);
  gl_rom_g35384 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_709(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_707(0), ZN => gl_rom_n_1036);
  gl_rom_g35385 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_1020(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_1018(1), ZN => gl_rom_n_1035);
  gl_rom_g35386 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_362(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_367(0), ZN => gl_rom_n_1034);
  gl_rom_g35387 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_704(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_705(0), ZN => gl_rom_n_1033);
  gl_rom_g35388 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_1017(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_1021(1), ZN => gl_rom_n_1032);
  gl_rom_g35389 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_1016(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_1019(1), ZN => gl_rom_n_1031);
  gl_rom_g35390 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_361(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_365(0), ZN => gl_rom_n_1030);
  gl_rom_g35391 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_1006(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_1007(1), ZN => gl_rom_n_1029);
  gl_rom_g35392 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_997(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_995(0), ZN => gl_rom_n_1028);
  gl_rom_g35393 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_1004(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_1002(1), ZN => gl_rom_n_1027);
  gl_rom_g35394 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_364(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_366(0), ZN => gl_rom_n_1026);
  gl_rom_g35395 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_360(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_363(0), ZN => gl_rom_n_1025);
  gl_rom_g35396 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_1001(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_1005(1), ZN => gl_rom_n_1024);
  gl_rom_g35397 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_1000(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_1003(1), ZN => gl_rom_n_1023);
  gl_rom_g35398 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_974(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_975(1), ZN => gl_rom_n_1022);
  gl_rom_g35399 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_957(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_955(0), ZN => gl_rom_n_1021);
  gl_rom_g35400 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_972(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_970(1), ZN => gl_rom_n_1020);
  gl_rom_g35401 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_370(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_375(0), ZN => gl_rom_n_1019);
  gl_rom_g35402 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_969(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_973(1), ZN => gl_rom_n_1018);
  gl_rom_g35403 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_854(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_855(0), ZN => gl_rom_n_1017);
  gl_rom_g35404 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_968(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_971(1), ZN => gl_rom_n_1016);
  gl_rom_g35405 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_372(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_374(0), ZN => gl_rom_n_1015);
  gl_rom_g35406 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_794(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_799(0), ZN => gl_rom_n_1014);
  gl_rom_g35407 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_966(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_967(1), ZN => gl_rom_n_1013);
  gl_rom_g35408 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_373(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_371(0), ZN => gl_rom_n_1012);
  gl_rom_g35409 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_964(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_962(1), ZN => gl_rom_n_1011);
  gl_rom_g35410 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_852(0), B1 => gl_rom_n_20, B2 => gl_rom_rom_850(0), ZN => gl_rom_n_1010);
  gl_rom_g35411 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_961(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_965(1), ZN => gl_rom_n_1009);
  gl_rom_g35412 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_960(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_963(1), ZN => gl_rom_n_1008);
  gl_rom_g35413 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_368(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_369(0), ZN => gl_rom_n_1007);
  gl_rom_g35414 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_953(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_957(1), ZN => gl_rom_n_1006);
  gl_rom_g35415 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_793(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_797(0), ZN => gl_rom_n_1005);
  gl_rom_g35416 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_796(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_798(0), ZN => gl_rom_n_1004);
  gl_rom_g35417 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_956(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_958(1), ZN => gl_rom_n_1003);
  gl_rom_g35418 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_338(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_343(0), ZN => gl_rom_n_1002);
  gl_rom_g35419 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_954(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_955(1), ZN => gl_rom_n_1001);
  gl_rom_g35420 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_340(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_342(0), ZN => gl_rom_n_1000);
  gl_rom_g35421 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_952(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_959(1), ZN => gl_rom_n_999);
  gl_rom_g35422 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_792(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_795(0), ZN => gl_rom_n_998);
  gl_rom_g35423 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_937(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_941(1), ZN => gl_rom_n_997);
  gl_rom_g35424 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_341(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_339(0), ZN => gl_rom_n_996);
  gl_rom_g35425 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_940(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_942(1), ZN => gl_rom_n_995);
  gl_rom_g35426 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_938(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_939(1), ZN => gl_rom_n_994);
  gl_rom_g35427 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_336(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_337(0), ZN => gl_rom_n_993);
  gl_rom_g35428 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_936(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_943(1), ZN => gl_rom_n_992);
  gl_rom_g35429 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_926(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_927(1), ZN => gl_rom_n_991);
  gl_rom_g35430 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_849(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_853(0), ZN => gl_rom_n_990);
  gl_rom_g35431 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_924(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_922(1), ZN => gl_rom_n_989);
  gl_rom_g35432 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_952(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_953(0), ZN => gl_rom_n_988);
  gl_rom_g35433 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_346(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_351(0), ZN => gl_rom_n_987);
  gl_rom_g35434 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_921(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_925(1), ZN => gl_rom_n_986);
  gl_rom_g35435 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_801(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_805(0), ZN => gl_rom_n_985);
  gl_rom_g35436 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_920(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_923(1), ZN => gl_rom_n_984);
  gl_rom_g35437 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_348(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_350(0), ZN => gl_rom_n_983);
  gl_rom_g35438 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_848(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_851(0), ZN => gl_rom_n_982);
  gl_rom_g35439 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_930(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_935(1), ZN => gl_rom_n_981);
  gl_rom_g35440 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_929(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_933(1), ZN => gl_rom_n_980);
  gl_rom_g35441 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_349(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_347(0), ZN => gl_rom_n_979);
  gl_rom_g35442 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_932(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_934(1), ZN => gl_rom_n_978);
  gl_rom_g35443 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_344(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_345(0), ZN => gl_rom_n_977);
  gl_rom_g35444 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_928(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_931(1), ZN => gl_rom_n_976);
  gl_rom_g35445 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_804(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_806(0), ZN => gl_rom_n_975);
  gl_rom_g35446 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_945(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_949(1), ZN => gl_rom_n_974);
  gl_rom_g35447 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_992(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_993(0), ZN => gl_rom_n_973);
  gl_rom_g35448 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_948(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_950(1), ZN => gl_rom_n_972);
  gl_rom_g35449 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_354(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_359(0), ZN => gl_rom_n_971);
  gl_rom_g35450 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_802(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_807(0), ZN => gl_rom_n_970);
  gl_rom_g35451 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_946(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_947(1), ZN => gl_rom_n_969);
  gl_rom_g35452 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_356(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_358(0), ZN => gl_rom_n_968);
  gl_rom_g35453 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_944(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_951(1), ZN => gl_rom_n_967);
  gl_rom_g35454 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_914(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_919(1), ZN => gl_rom_n_966);
  gl_rom_g35455 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_800(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_803(0), ZN => gl_rom_n_965);
  gl_rom_g35456 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_357(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_355(0), ZN => gl_rom_n_964);
  gl_rom_g35457 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_913(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_917(1), ZN => gl_rom_n_963);
  gl_rom_g35458 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_352(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_353(0), ZN => gl_rom_n_962);
  gl_rom_g35459 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_916(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_915(1), ZN => gl_rom_n_961);
  gl_rom_g35460 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_912(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_918(1), ZN => gl_rom_n_960);
  gl_rom_g35461 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_905(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_909(1), ZN => gl_rom_n_959);
  gl_rom_g35462 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_908(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_910(1), ZN => gl_rom_n_958);
  gl_rom_g35463 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_329(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_333(0), ZN => gl_rom_n_957);
  gl_rom_g35464 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_906(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_911(1), ZN => gl_rom_n_956);
  gl_rom_g35465 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_904(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_907(1), ZN => gl_rom_n_955);
  gl_rom_g35466 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_332(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_334(0), ZN => gl_rom_n_954);
  gl_rom_g35467 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_817(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_821(0), ZN => gl_rom_n_953);
  gl_rom_g35468 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_938(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_943(0), ZN => gl_rom_n_952);
  gl_rom_g35469 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_898(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_903(1), ZN => gl_rom_n_951);
  gl_rom_g35470 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_890(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_895(0), ZN => gl_rom_n_950);
  gl_rom_g35471 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_330(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_331(0), ZN => gl_rom_n_949);
  gl_rom_g35472 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_897(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_901(1), ZN => gl_rom_n_948);
  gl_rom_g35473 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_820(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_822(0), ZN => gl_rom_n_947);
  gl_rom_g35474 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_328(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_335(0), ZN => gl_rom_n_946);
  gl_rom_g35475 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_900(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_902(1), ZN => gl_rom_n_945);
  gl_rom_g35476 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_896(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_899(1), ZN => gl_rom_n_944);
  gl_rom_g35477 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_892(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_894(0), ZN => gl_rom_n_943);
  gl_rom_g35478 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_702(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_703(1), ZN => gl_rom_n_942);
  gl_rom_g35479 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_322(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_327(0), ZN => gl_rom_n_941);
  gl_rom_g35480 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_700(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_698(1), ZN => gl_rom_n_940);
  gl_rom_g35481 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_818(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_819(0), ZN => gl_rom_n_939);
  gl_rom_g35482 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_697(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_701(1), ZN => gl_rom_n_938);
  gl_rom_g35483 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_696(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_699(1), ZN => gl_rom_n_937);
  gl_rom_g35484 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_324(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_326(0), ZN => gl_rom_n_936);
  gl_rom_g35485 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_325(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_323(0), ZN => gl_rom_n_935);
  gl_rom_g35486 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_686(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_687(1), ZN => gl_rom_n_934);
  gl_rom_g35487 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_816(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_823(0), ZN => gl_rom_n_933);
  gl_rom_g35488 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_684(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_682(1), ZN => gl_rom_n_932);
  gl_rom_g35489 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_320(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_321(0), ZN => gl_rom_n_931);
  gl_rom_g35490 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_681(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_685(1), ZN => gl_rom_n_930);
  gl_rom_g35491 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_680(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_683(1), ZN => gl_rom_n_929);
  gl_rom_g35492 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_893(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_891(0), ZN => gl_rom_n_928);
  gl_rom_g35493 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_690(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_695(1), ZN => gl_rom_n_927);
  gl_rom_g35494 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_692(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_694(1), ZN => gl_rom_n_926);
  gl_rom_g35495 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_940(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_942(0), ZN => gl_rom_n_925);
  gl_rom_g35496 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_126(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_127(0), ZN => gl_rom_n_924);
  gl_rom_g35497 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_693(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_691(1), ZN => gl_rom_n_923);
  gl_rom_g35498 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_688(1), B1 => gl_rom_n_21, B2 => gl_rom_rom_689(1), ZN => gl_rom_n_922);
  gl_rom_g35499 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_124(0), B1 => gl_rom_n_20, B2 => gl_rom_rom_122(0), ZN => gl_rom_n_921);
  gl_rom_g35500 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_662(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_663(1), ZN => gl_rom_n_920);
  gl_rom_g35501 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_786(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_791(0), ZN => gl_rom_n_919);
  gl_rom_g35502 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_660(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_658(1), ZN => gl_rom_n_918);
  gl_rom_g35503 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_785(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_789(0), ZN => gl_rom_n_917);
  gl_rom_g35504 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_121(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_125(0), ZN => gl_rom_n_916);
  gl_rom_g35505 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_120(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_123(0), ZN => gl_rom_n_915);
  gl_rom_g35506 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_657(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_661(1), ZN => gl_rom_n_914);
  gl_rom_g35507 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_656(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_659(1), ZN => gl_rom_n_913);
  gl_rom_g35508 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_666(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_671(1), ZN => gl_rom_n_912);
  gl_rom_g35509 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_978(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_983(0), ZN => gl_rom_n_911);
  gl_rom_g35510 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_888(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_889(0), ZN => gl_rom_n_910);
  gl_rom_g35511 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_788(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_787(0), ZN => gl_rom_n_909);
  gl_rom_g35512 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_665(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_669(1), ZN => gl_rom_n_908);
  gl_rom_g35513 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_106(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_111(0), ZN => gl_rom_n_907);
  gl_rom_g35514 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_105(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_109(0), ZN => gl_rom_n_906);
  gl_rom_g35515 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_668(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_667(1), ZN => gl_rom_n_905);
  gl_rom_g35516 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_664(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_670(1), ZN => gl_rom_n_904);
  gl_rom_g35517 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_678(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_679(1), ZN => gl_rom_n_903);
  gl_rom_g35518 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_941(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_939(0), ZN => gl_rom_n_902);
  gl_rom_g35519 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_784(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_790(0), ZN => gl_rom_n_901);
  gl_rom_g35520 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_108(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_107(0), ZN => gl_rom_n_900);
  gl_rom_g35521 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_676(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_674(1), ZN => gl_rom_n_899);
  gl_rom_g35522 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_104(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_110(0), ZN => gl_rom_n_898);
  gl_rom_g35523 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_673(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_677(1), ZN => gl_rom_n_897);
  gl_rom_g35524 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_672(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_675(1), ZN => gl_rom_n_896);
  gl_rom_g35525 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_654(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_655(1), ZN => gl_rom_n_895);
  gl_rom_g35526 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_652(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_650(1), ZN => gl_rom_n_894);
  gl_rom_g35527 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_874(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_879(0), ZN => gl_rom_n_893);
  gl_rom_g35528 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_114(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_119(0), ZN => gl_rom_n_892);
  gl_rom_g35529 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_649(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_653(1), ZN => gl_rom_n_891);
  gl_rom_g35530 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_116(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_118(0), ZN => gl_rom_n_890);
  gl_rom_g35531 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_648(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_651(1), ZN => gl_rom_n_889);
  gl_rom_g35532 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_825(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_829(0), ZN => gl_rom_n_888);
  gl_rom_g35533 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_828(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_830(0), ZN => gl_rom_n_887);
  gl_rom_g35534 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_642(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_647(1), ZN => gl_rom_n_886);
  gl_rom_g35535 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_117(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_115(0), ZN => gl_rom_n_885);
  gl_rom_g35536 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_641(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_645(1), ZN => gl_rom_n_884);
  gl_rom_g35537 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_644(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_646(1), ZN => gl_rom_n_883);
  gl_rom_g35538 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_640(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_643(1), ZN => gl_rom_n_882);
  gl_rom_g35539 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_569(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_573(1), ZN => gl_rom_n_881);
  gl_rom_g35540 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_112(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_113(0), ZN => gl_rom_n_880);
  gl_rom_g35541 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_873(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_877(0), ZN => gl_rom_n_879);
  gl_rom_g35542 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_82(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_87(0), ZN => gl_rom_n_878);
  gl_rom_g35543 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_572(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_574(1), ZN => gl_rom_n_877);
  gl_rom_g35544 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_826(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_827(0), ZN => gl_rom_n_876);
  gl_rom_g35545 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_570(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_571(1), ZN => gl_rom_n_875);
  gl_rom_g35546 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_84(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_86(0), ZN => gl_rom_n_874);
  gl_rom_g35547 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_568(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_575(1), ZN => gl_rom_n_873);
  gl_rom_g35548 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_824(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_831(0), ZN => gl_rom_n_872);
  gl_rom_g35549 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_85(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_83(0), ZN => gl_rom_n_871);
  gl_rom_g35550 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_554(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_559(1), ZN => gl_rom_n_870);
  gl_rom_g35551 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_553(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_557(1), ZN => gl_rom_n_869);
  gl_rom_g35552 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_556(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_558(1), ZN => gl_rom_n_868);
  gl_rom_g35553 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_80(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_81(0), ZN => gl_rom_n_867);
  gl_rom_g35554 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_552(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_555(1), ZN => gl_rom_n_866);
  gl_rom_g35555 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_936(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_937(0), ZN => gl_rom_n_865);
  gl_rom_g35556 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_876(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_875(0), ZN => gl_rom_n_864);
  gl_rom_g35557 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_566(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_567(1), ZN => gl_rom_n_863);
  gl_rom_g35558 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_980(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_982(0), ZN => gl_rom_n_862);
  gl_rom_g35559 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_1018(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_1023(0), ZN => gl_rom_n_861);
  gl_rom_g35560 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_564(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_562(1), ZN => gl_rom_n_860);
  gl_rom_g35561 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_90(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_95(0), ZN => gl_rom_n_859);
  gl_rom_g35562 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_810(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_815(0), ZN => gl_rom_n_858);
  gl_rom_g35563 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_561(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_565(1), ZN => gl_rom_n_857);
  gl_rom_g35564 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_92(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_94(0), ZN => gl_rom_n_856);
  gl_rom_g35565 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_560(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_563(1), ZN => gl_rom_n_855);
  gl_rom_g35566 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_534(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_535(1), ZN => gl_rom_n_854);
  gl_rom_g35567 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_93(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_91(0), ZN => gl_rom_n_853);
  gl_rom_g35568 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_532(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_530(1), ZN => gl_rom_n_852);
  gl_rom_g35569 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_809(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_813(0), ZN => gl_rom_n_851);
  gl_rom_g35570 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_529(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_533(1), ZN => gl_rom_n_850);
  gl_rom_g35571 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_528(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_531(1), ZN => gl_rom_n_849);
  gl_rom_g35572 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_88(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_89(0), ZN => gl_rom_n_848);
  gl_rom_g35573 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_542(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_543(1), ZN => gl_rom_n_847);
  gl_rom_g35574 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_872(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_878(0), ZN => gl_rom_n_846);
  gl_rom_g35575 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_812(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_811(0), ZN => gl_rom_n_845);
  gl_rom_g35576 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_102(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_103(0), ZN => gl_rom_n_844);
  gl_rom_g35577 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_540(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_538(1), ZN => gl_rom_n_843);
  gl_rom_g35578 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_100(0), B1 => gl_rom_n_20, B2 => gl_rom_rom_98(0), ZN => gl_rom_n_842);
  gl_rom_g35579 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_537(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_541(1), ZN => gl_rom_n_841);
  gl_rom_g35580 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_536(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_539(1), ZN => gl_rom_n_840);
  gl_rom_g35581 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_550(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_551(1), ZN => gl_rom_n_839);
  gl_rom_g35582 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_808(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_814(0), ZN => gl_rom_n_838);
  gl_rom_g35583 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_97(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_101(0), ZN => gl_rom_n_837);
  gl_rom_g35584 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_548(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_546(1), ZN => gl_rom_n_836);
  gl_rom_g35585 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_96(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_99(0), ZN => gl_rom_n_835);
  gl_rom_g35586 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_545(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_549(1), ZN => gl_rom_n_834);
  gl_rom_g35587 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_544(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_547(1), ZN => gl_rom_n_833);
  gl_rom_g35588 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_526(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_527(1), ZN => gl_rom_n_832);
  gl_rom_g35589 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_524(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_522(1), ZN => gl_rom_n_831);
  gl_rom_g35590 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_74(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_79(0), ZN => gl_rom_n_830);
  gl_rom_g35591 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_842(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_847(0), ZN => gl_rom_n_829);
  gl_rom_g35592 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_521(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_525(1), ZN => gl_rom_n_828);
  gl_rom_g35593 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_778(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_783(0), ZN => gl_rom_n_827);
  gl_rom_g35594 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_520(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_523(1), ZN => gl_rom_n_826);
  gl_rom_g35595 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_73(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_77(0), ZN => gl_rom_n_825);
  gl_rom_g35596 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_946(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_951(0), ZN => gl_rom_n_824);
  gl_rom_g35597 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_513(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_517(1), ZN => gl_rom_n_823);
  gl_rom_g35598 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_76(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_75(0), ZN => gl_rom_n_822);
  gl_rom_g35599 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_516(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_518(1), ZN => gl_rom_n_821);
  gl_rom_g35600 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_72(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_78(0), ZN => gl_rom_n_820);
  gl_rom_g35601 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_514(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_519(1), ZN => gl_rom_n_819);
  gl_rom_g35602 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_512(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_515(1), ZN => gl_rom_n_818);
  gl_rom_g35603 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_777(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_781(0), ZN => gl_rom_n_817);
  gl_rom_g35604 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_1017(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_1021(0), ZN => gl_rom_n_816);
  gl_rom_g35605 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_66(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_71(0), ZN => gl_rom_n_815);
  gl_rom_g35606 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_780(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_782(0), ZN => gl_rom_n_814);
  gl_rom_g35607 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_498(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_503(1), ZN => gl_rom_n_813);
  gl_rom_g35608 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_497(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_501(1), ZN => gl_rom_n_812);
  gl_rom_g35609 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_841(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_845(0), ZN => gl_rom_n_811);
  gl_rom_g35610 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_68(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_70(0), ZN => gl_rom_n_810);
  gl_rom_g35611 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_500(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_502(1), ZN => gl_rom_n_809);
  gl_rom_g35612 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_496(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_499(1), ZN => gl_rom_n_808);
  gl_rom_g35613 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_69(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_67(0), ZN => gl_rom_n_807);
  gl_rom_g35614 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_1008(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_1011(1), ZN => gl_rom_n_806);
  gl_rom_g35615 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_465(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_469(1), ZN => gl_rom_n_805);
  gl_rom_g35616 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_468(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_470(1), ZN => gl_rom_n_804);
  gl_rom_g35617 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_64(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_65(0), ZN => gl_rom_n_803);
  gl_rom_g35618 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_466(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_471(1), ZN => gl_rom_n_802);
  gl_rom_g35619 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_464(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_467(1), ZN => gl_rom_n_801);
  gl_rom_g35620 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_844(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_843(0), ZN => gl_rom_n_800);
  gl_rom_g35621 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_474(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_479(1), ZN => gl_rom_n_799);
  gl_rom_g35622 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_945(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_949(0), ZN => gl_rom_n_798);
  gl_rom_g35623 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_770(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_775(0), ZN => gl_rom_n_797);
  gl_rom_g35624 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_476(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_478(1), ZN => gl_rom_n_796);
  gl_rom_g35625 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_217(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_221(0), ZN => gl_rom_n_795);
  gl_rom_g35626 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_477(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_475(1), ZN => gl_rom_n_794);
  gl_rom_g35627 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_472(1), B1 => gl_rom_n_21, B2 => gl_rom_rom_473(1), ZN => gl_rom_n_793);
  gl_rom_g35628 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_220(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_222(0), ZN => gl_rom_n_792);
  gl_rom_g35629 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_769(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_773(0), ZN => gl_rom_n_791);
  gl_rom_g35630 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_486(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_487(1), ZN => gl_rom_n_790);
  gl_rom_g35631 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_484(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_482(1), ZN => gl_rom_n_789);
  gl_rom_g35632 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_218(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_219(0), ZN => gl_rom_n_788);
  gl_rom_g35633 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_481(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_485(1), ZN => gl_rom_n_787);
  gl_rom_g35634 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_480(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_483(1), ZN => gl_rom_n_786);
  gl_rom_g35635 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_216(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_223(0), ZN => gl_rom_n_785);
  gl_rom_g35636 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_506(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_511(1), ZN => gl_rom_n_784);
  gl_rom_g35637 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_840(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_846(0), ZN => gl_rom_n_783);
  gl_rom_g35638 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_772(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_774(0), ZN => gl_rom_n_782);
  gl_rom_g35639 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_225(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_229(0), ZN => gl_rom_n_781);
  gl_rom_g35640 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_508(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_510(1), ZN => gl_rom_n_780);
  gl_rom_g35641 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_768(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_771(0), ZN => gl_rom_n_779);
  gl_rom_g35642 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_509(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_507(1), ZN => gl_rom_n_778);
  gl_rom_g35643 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_228(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_230(0), ZN => gl_rom_n_777);
  gl_rom_g35644 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_504(1), B1 => gl_rom_n_21, B2 => gl_rom_rom_505(1), ZN => gl_rom_n_776);
  gl_rom_g35645 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_489(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_493(1), ZN => gl_rom_n_775);
  gl_rom_g35646 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_226(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_227(0), ZN => gl_rom_n_774);
  gl_rom_g35647 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_492(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_494(1), ZN => gl_rom_n_773);
  gl_rom_g35648 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_1012(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_1014(0), ZN => gl_rom_n_772);
  gl_rom_g35649 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_490(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_495(1), ZN => gl_rom_n_771);
  gl_rom_g35650 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_224(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_231(0), ZN => gl_rom_n_770);
  gl_rom_g35651 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_488(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_491(1), ZN => gl_rom_n_769);
  gl_rom_g35652 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_948(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_947(0), ZN => gl_rom_n_768);
  gl_rom_g35653 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_834(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_839(0), ZN => gl_rom_n_767);
  gl_rom_g35654 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_458(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_463(1), ZN => gl_rom_n_766);
  gl_rom_g35655 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_457(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_461(1), ZN => gl_rom_n_765);
  gl_rom_g35656 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_242(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_247(0), ZN => gl_rom_n_764);
  gl_rom_g35657 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_460(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_462(1), ZN => gl_rom_n_763);
  gl_rom_g35658 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_456(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_459(1), ZN => gl_rom_n_762);
  gl_rom_g35659 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_241(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_245(0), ZN => gl_rom_n_761);
  gl_rom_g35660 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_702(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_703(0), ZN => gl_rom_n_760);
  gl_rom_g35661 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_449(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_453(1), ZN => gl_rom_n_759);
  gl_rom_g35662 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_244(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_246(0), ZN => gl_rom_n_758);
  gl_rom_g35663 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_452(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_454(1), ZN => gl_rom_n_757);
  gl_rom_g35664 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_981(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_979(0), ZN => gl_rom_n_756);
  gl_rom_g35665 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_450(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_455(1), ZN => gl_rom_n_755);
  gl_rom_g35666 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_240(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_243(0), ZN => gl_rom_n_754);
  gl_rom_g35667 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_448(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_451(1), ZN => gl_rom_n_753);
  gl_rom_g35668 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_833(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_837(0), ZN => gl_rom_n_752);
  gl_rom_g35669 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_700(0), B1 => gl_rom_n_20, B2 => gl_rom_rom_698(0), ZN => gl_rom_n_751);
  gl_rom_g35670 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_442(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_447(1), ZN => gl_rom_n_750);
  gl_rom_g35671 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_214(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_215(0), ZN => gl_rom_n_749);
  gl_rom_g35672 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_444(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_446(1), ZN => gl_rom_n_748);
  gl_rom_g35673 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_212(0), B1 => gl_rom_n_20, B2 => gl_rom_rom_210(0), ZN => gl_rom_n_747);
  gl_rom_g35674 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_445(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_443(1), ZN => gl_rom_n_746);
  gl_rom_g35675 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_440(1), B1 => gl_rom_n_21, B2 => gl_rom_rom_441(1), ZN => gl_rom_n_745);
  gl_rom_g35676 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_697(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_701(0), ZN => gl_rom_n_744);
  gl_rom_g35677 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_1020(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_1022(0), ZN => gl_rom_n_743);
  gl_rom_g35678 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_944(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_950(0), ZN => gl_rom_n_742);
  gl_rom_g35679 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_426(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_431(1), ZN => gl_rom_n_741);
  gl_rom_g35680 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_209(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_213(0), ZN => gl_rom_n_740);
  gl_rom_g35681 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_425(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_429(1), ZN => gl_rom_n_739);
  gl_rom_g35682 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_428(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_430(1), ZN => gl_rom_n_738);
  gl_rom_g35683 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_424(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_427(1), ZN => gl_rom_n_737);
  gl_rom_g35684 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_208(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_211(0), ZN => gl_rom_n_736);
  gl_rom_g35685 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_836(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_835(0), ZN => gl_rom_n_735);
  gl_rom_g35686 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_410(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_415(1), ZN => gl_rom_n_734);
  gl_rom_g35687 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_409(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_413(1), ZN => gl_rom_n_733);
  gl_rom_g35688 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_696(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_699(0), ZN => gl_rom_n_732);
  gl_rom_g35689 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_254(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_255(0), ZN => gl_rom_n_731);
  gl_rom_g35690 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_412(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_414(1), ZN => gl_rom_n_730);
  gl_rom_g35691 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_252(0), B1 => gl_rom_n_20, B2 => gl_rom_rom_250(0), ZN => gl_rom_n_729);
  gl_rom_g35692 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_408(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_411(1), ZN => gl_rom_n_728);
  gl_rom_g35693 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_681(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_685(0), ZN => gl_rom_n_727);
  gl_rom_g35694 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_832(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_838(0), ZN => gl_rom_n_726);
  gl_rom_g35695 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_422(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_423(1), ZN => gl_rom_n_725);
  gl_rom_g35696 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_249(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_253(0), ZN => gl_rom_n_724);
  gl_rom_g35697 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_420(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_418(1), ZN => gl_rom_n_723);
  gl_rom_g35698 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_684(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_686(0), ZN => gl_rom_n_722);
  gl_rom_g35699 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_417(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_421(1), ZN => gl_rom_n_721);
  gl_rom_g35700 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_416(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_419(1), ZN => gl_rom_n_720);
  gl_rom_g35701 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_248(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_251(0), ZN => gl_rom_n_719);
  gl_rom_g35702 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_433(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_437(1), ZN => gl_rom_n_718);
  gl_rom_g35703 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_436(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_438(1), ZN => gl_rom_n_717);
  gl_rom_g35704 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_233(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_237(0), ZN => gl_rom_n_716);
  gl_rom_g35705 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_434(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_439(1), ZN => gl_rom_n_715);
  gl_rom_g35706 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_236(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_238(0), ZN => gl_rom_n_714);
  gl_rom_g35707 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_432(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_435(1), ZN => gl_rom_n_713);
  gl_rom_g35708 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_682(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_683(0), ZN => gl_rom_n_712);
  gl_rom_g35709 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_402(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_407(1), ZN => gl_rom_n_711);
  gl_rom_g35710 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_234(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_235(0), ZN => gl_rom_n_710);
  gl_rom_g35711 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_401(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_405(1), ZN => gl_rom_n_709);
  gl_rom_g35712 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_680(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_687(0), ZN => gl_rom_n_708);
  gl_rom_g35713 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_404(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_406(1), ZN => gl_rom_n_707);
  gl_rom_g35714 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_1016(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_1019(0), ZN => gl_rom_n_706);
  gl_rom_g35715 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_232(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_239(0), ZN => gl_rom_n_705);
  gl_rom_g35716 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_400(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_403(1), ZN => gl_rom_n_704);
  gl_rom_g35717 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_914(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_919(0), ZN => gl_rom_n_703);
  gl_rom_g35718 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_393(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_397(1), ZN => gl_rom_n_702);
  gl_rom_g35719 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_396(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_398(1), ZN => gl_rom_n_701);
  gl_rom_g35720 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_201(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_205(0), ZN => gl_rom_n_700);
  gl_rom_g35721 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_394(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_399(1), ZN => gl_rom_n_699);
  gl_rom_g35722 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_916(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_918(0), ZN => gl_rom_n_698);
  gl_rom_g35723 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_204(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_206(0), ZN => gl_rom_n_697);
  gl_rom_g35724 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_392(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_395(1), ZN => gl_rom_n_696);
  gl_rom_g35725 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_666(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_671(0), ZN => gl_rom_n_695);
  gl_rom_g35726 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_390(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_391(1), ZN => gl_rom_n_694);
  gl_rom_g35727 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_634(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_639(0), ZN => gl_rom_n_693);
  gl_rom_g35728 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_388(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_386(1), ZN => gl_rom_n_692);
  gl_rom_g35729 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_202(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_203(0), ZN => gl_rom_n_691);
  gl_rom_g35730 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_385(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_389(1), ZN => gl_rom_n_690);
  gl_rom_g35731 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_668(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_670(0), ZN => gl_rom_n_689);
  gl_rom_g35732 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_200(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_207(0), ZN => gl_rom_n_688);
  gl_rom_g35733 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_384(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_387(1), ZN => gl_rom_n_687);
  gl_rom_g35734 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_193(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_197(0), ZN => gl_rom_n_686);
  gl_rom_g35735 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_249(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_253(1), ZN => gl_rom_n_685);
  gl_rom_g35736 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_252(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_254(1), ZN => gl_rom_n_684);
  gl_rom_g35737 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_669(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_667(0), ZN => gl_rom_n_683);
  gl_rom_g35738 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_196(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_198(0), ZN => gl_rom_n_682);
  gl_rom_g35739 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_250(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_251(1), ZN => gl_rom_n_681);
  gl_rom_g35740 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_248(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_255(1), ZN => gl_rom_n_680);
  gl_rom_g35741 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_636(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_638(0), ZN => gl_rom_n_679);
  gl_rom_g35742 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_194(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_195(0), ZN => gl_rom_n_678);
  gl_rom_g35743 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_234(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_239(1), ZN => gl_rom_n_677);
  gl_rom_g35744 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_233(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_237(1), ZN => gl_rom_n_676);
  gl_rom_g35745 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_192(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_199(0), ZN => gl_rom_n_675);
  gl_rom_g35746 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_236(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_235(1), ZN => gl_rom_n_674);
  gl_rom_g35747 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_232(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_238(1), ZN => gl_rom_n_673);
  gl_rom_g35748 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_664(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_665(0), ZN => gl_rom_n_672);
  gl_rom_g35749 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_241(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_245(1), ZN => gl_rom_n_671);
  gl_rom_g35750 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_244(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_246(1), ZN => gl_rom_n_670);
  gl_rom_g35751 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_637(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_635(0), ZN => gl_rom_n_669);
  gl_rom_g35752 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_318(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_319(0), ZN => gl_rom_n_668);
  gl_rom_g35753 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_242(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_243(1), ZN => gl_rom_n_667);
  gl_rom_g35754 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_240(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_247(1), ZN => gl_rom_n_666);
  gl_rom_g35755 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_674(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_679(0), ZN => gl_rom_n_665);
  gl_rom_g35756 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_316(0), B1 => gl_rom_n_20, B2 => gl_rom_rom_314(0), ZN => gl_rom_n_664);
  gl_rom_g35757 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_676(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_678(0), ZN => gl_rom_n_663);
  gl_rom_g35758 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_214(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_215(1), ZN => gl_rom_n_662);
  gl_rom_g35759 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_212(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_210(1), ZN => gl_rom_n_661);
  gl_rom_g35760 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_313(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_317(0), ZN => gl_rom_n_660);
  gl_rom_g35761 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_209(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_213(1), ZN => gl_rom_n_659);
  gl_rom_g35762 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_208(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_211(1), ZN => gl_rom_n_658);
  gl_rom_g35763 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_312(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_315(0), ZN => gl_rom_n_657);
  gl_rom_g35764 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_218(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_223(1), ZN => gl_rom_n_656);
  gl_rom_g35765 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_677(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_675(0), ZN => gl_rom_n_655);
  gl_rom_g35766 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_217(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_221(1), ZN => gl_rom_n_654);
  gl_rom_g35767 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_302(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_303(0), ZN => gl_rom_n_653);
  gl_rom_g35768 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_632(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_633(0), ZN => gl_rom_n_652);
  gl_rom_g35769 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_220(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_222(1), ZN => gl_rom_n_651);
  gl_rom_g35770 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_300(0), B1 => gl_rom_n_20, B2 => gl_rom_rom_298(0), ZN => gl_rom_n_650);
  gl_rom_g35771 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_216(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_219(1), ZN => gl_rom_n_649);
  gl_rom_g35772 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_672(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_673(0), ZN => gl_rom_n_648);
  gl_rom_g35773 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_226(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_231(1), ZN => gl_rom_n_647);
  gl_rom_g35774 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_228(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_230(1), ZN => gl_rom_n_646);
  gl_rom_g35775 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_297(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_301(0), ZN => gl_rom_n_645);
  gl_rom_g35776 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_229(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_227(1), ZN => gl_rom_n_644);
  gl_rom_g35777 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_296(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_299(0), ZN => gl_rom_n_643);
  gl_rom_g35778 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_224(1), B1 => gl_rom_n_21, B2 => gl_rom_rom_225(1), ZN => gl_rom_n_642);
  gl_rom_g35779 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_976(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_977(0), ZN => gl_rom_n_641);
  gl_rom_g35780 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_202(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_207(1), ZN => gl_rom_n_640);
  gl_rom_g35781 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_917(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_915(0), ZN => gl_rom_n_639);
  gl_rom_g35782 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_201(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_205(1), ZN => gl_rom_n_638);
  gl_rom_g35783 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_281(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_285(0), ZN => gl_rom_n_637);
  gl_rom_g35784 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_912(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_913(0), ZN => gl_rom_n_636);
  gl_rom_g35785 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_204(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_206(1), ZN => gl_rom_n_635);
  gl_rom_g35786 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_200(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_203(1), ZN => gl_rom_n_634);
  gl_rom_g35787 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_284(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_286(0), ZN => gl_rom_n_633);
  gl_rom_g35788 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_689(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_693(0), ZN => gl_rom_n_632);
  gl_rom_g35789 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_193(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_197(1), ZN => gl_rom_n_631);
  gl_rom_g35790 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_282(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_283(0), ZN => gl_rom_n_630);
  gl_rom_g35791 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_196(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_198(1), ZN => gl_rom_n_629);
  gl_rom_g35792 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_617(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_621(0), ZN => gl_rom_n_628);
  gl_rom_g35793 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_280(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_287(0), ZN => gl_rom_n_627);
  gl_rom_g35794 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_194(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_195(1), ZN => gl_rom_n_626);
  gl_rom_g35795 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_192(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_199(1), ZN => gl_rom_n_625);
  gl_rom_g35796 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_692(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_694(0), ZN => gl_rom_n_624);
  gl_rom_g35797 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_620(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_622(0), ZN => gl_rom_n_623);
  gl_rom_g35798 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_318(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_319(1), ZN => gl_rom_n_622);
  gl_rom_g35799 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_289(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_293(0), ZN => gl_rom_n_621);
  gl_rom_g35800 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_316(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_314(1), ZN => gl_rom_n_620);
  gl_rom_g35801 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_690(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_695(0), ZN => gl_rom_n_619);
  gl_rom_g35802 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_292(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_294(0), ZN => gl_rom_n_618);
  gl_rom_g35803 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_313(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_317(1), ZN => gl_rom_n_617);
  gl_rom_g35804 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_688(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_691(0), ZN => gl_rom_n_616);
  gl_rom_g35805 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_312(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_315(1), ZN => gl_rom_n_615);
  gl_rom_g35806 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_290(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_291(0), ZN => gl_rom_n_614);
  gl_rom_g35807 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_302(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_303(1), ZN => gl_rom_n_613);
  gl_rom_g35808 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_300(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_298(1), ZN => gl_rom_n_612);
  gl_rom_g35809 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_297(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_301(1), ZN => gl_rom_n_611);
  gl_rom_g35810 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_296(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_299(1), ZN => gl_rom_n_610);
  gl_rom_g35811 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_288(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_295(0), ZN => gl_rom_n_609);
  gl_rom_g35812 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_618(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_619(0), ZN => gl_rom_n_608);
  gl_rom_g35813 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_310(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_311(1), ZN => gl_rom_n_607);
  gl_rom_g35814 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_308(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_306(1), ZN => gl_rom_n_606);
  gl_rom_g35815 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_306(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_311(0), ZN => gl_rom_n_605);
  gl_rom_g35816 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_1001(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_1005(0), ZN => gl_rom_n_604);
  gl_rom_g35817 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_305(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_309(1), ZN => gl_rom_n_603);
  gl_rom_g35818 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_304(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_307(1), ZN => gl_rom_n_602);
  gl_rom_g35819 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_308(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_310(0), ZN => gl_rom_n_601);
  gl_rom_g35820 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_658(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_663(0), ZN => gl_rom_n_600);
  gl_rom_g35821 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_274(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_279(1), ZN => gl_rom_n_599);
  gl_rom_g35822 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_309(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_307(0), ZN => gl_rom_n_598);
  gl_rom_g35823 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_273(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_277(1), ZN => gl_rom_n_597);
  gl_rom_g35824 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_657(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_661(0), ZN => gl_rom_n_596);
  gl_rom_g35825 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_276(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_278(1), ZN => gl_rom_n_595);
  gl_rom_g35826 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_272(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_275(1), ZN => gl_rom_n_594);
  gl_rom_g35827 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_304(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_305(0), ZN => gl_rom_n_593);
  gl_rom_g35828 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_282(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_287(1), ZN => gl_rom_n_592);
  gl_rom_g35829 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_274(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_279(0), ZN => gl_rom_n_591);
  gl_rom_g35830 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_281(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_285(1), ZN => gl_rom_n_590);
  gl_rom_g35831 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_616(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_623(0), ZN => gl_rom_n_589);
  gl_rom_g35832 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_660(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_659(0), ZN => gl_rom_n_588);
  gl_rom_g35833 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_284(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_286(1), ZN => gl_rom_n_587);
  gl_rom_g35834 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_280(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_283(1), ZN => gl_rom_n_586);
  gl_rom_g35835 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_273(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_277(0), ZN => gl_rom_n_585);
  gl_rom_g35836 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_276(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_275(0), ZN => gl_rom_n_584);
  gl_rom_g35837 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_290(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_295(1), ZN => gl_rom_n_583);
  gl_rom_g35838 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_289(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_293(1), ZN => gl_rom_n_582);
  gl_rom_g35839 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_656(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_662(0), ZN => gl_rom_n_581);
  gl_rom_g35840 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_292(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_294(1), ZN => gl_rom_n_580);
  gl_rom_g35841 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_272(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_278(0), ZN => gl_rom_n_579);
  gl_rom_g35842 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_288(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_291(1), ZN => gl_rom_n_578);
  gl_rom_g35843 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_1004(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_1006(0), ZN => gl_rom_n_577);
  gl_rom_g35844 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_270(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_271(1), ZN => gl_rom_n_576);
  gl_rom_g35845 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_921(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_925(0), ZN => gl_rom_n_575);
  gl_rom_g35846 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_266(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_271(0), ZN => gl_rom_n_574);
  gl_rom_g35847 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_268(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_266(1), ZN => gl_rom_n_573);
  gl_rom_g35848 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_265(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_269(1), ZN => gl_rom_n_572);
  gl_rom_g35849 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_654(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_655(0), ZN => gl_rom_n_571);
  gl_rom_g35850 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_268(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_270(0), ZN => gl_rom_n_570);
  gl_rom_g35851 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_264(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_267(1), ZN => gl_rom_n_569);
  gl_rom_g35852 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_602(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_607(0), ZN => gl_rom_n_568);
  gl_rom_g35853 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_258(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_263(1), ZN => gl_rom_n_567);
  gl_rom_g35854 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_269(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_267(0), ZN => gl_rom_n_566);
  gl_rom_g35855 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_257(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_261(1), ZN => gl_rom_n_565);
  gl_rom_g35856 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_264(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_265(0), ZN => gl_rom_n_564);
  gl_rom_g35857 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_260(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_262(1), ZN => gl_rom_n_563);
  gl_rom_g35858 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_256(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_259(1), ZN => gl_rom_n_562);
  gl_rom_g35859 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_652(0), B1 => gl_rom_n_20, B2 => gl_rom_rom_650(0), ZN => gl_rom_n_561);
  gl_rom_g35860 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_258(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_263(0), ZN => gl_rom_n_560);
  gl_rom_g35861 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_346(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_351(1), ZN => gl_rom_n_559);
  gl_rom_g35862 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_604(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_606(0), ZN => gl_rom_n_558);
  gl_rom_g35863 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_345(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_349(1), ZN => gl_rom_n_557);
  gl_rom_g35864 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_257(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_261(0), ZN => gl_rom_n_556);
  gl_rom_g35865 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_348(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_350(1), ZN => gl_rom_n_555);
  gl_rom_g35866 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_649(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_653(0), ZN => gl_rom_n_554);
  gl_rom_g35867 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_344(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_347(1), ZN => gl_rom_n_553);
  gl_rom_g35868 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_260(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_259(0), ZN => gl_rom_n_552);
  gl_rom_g35869 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_648(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_651(0), ZN => gl_rom_n_551);
  gl_rom_g35870 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_892(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_890(1), ZN => gl_rom_n_550);
  gl_rom_g35871 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_356(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_358(1), ZN => gl_rom_n_549);
  gl_rom_g35872 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_256(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_262(0), ZN => gl_rom_n_548);
  gl_rom_g35873 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_354(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_355(1), ZN => gl_rom_n_547);
  gl_rom_g35874 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_352(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_359(1), ZN => gl_rom_n_546);
  gl_rom_g35875 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_924(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_926(0), ZN => gl_rom_n_545);
  gl_rom_g35876 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_370(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_375(1), ZN => gl_rom_n_544);
  gl_rom_g35877 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_369(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_373(1), ZN => gl_rom_n_543);
  gl_rom_g35878 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_605(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_603(0), ZN => gl_rom_n_542);
  gl_rom_g35879 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_190(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_191(0), ZN => gl_rom_n_541);
  gl_rom_g35880 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_641(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_645(0), ZN => gl_rom_n_540);
  gl_rom_g35881 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_372(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_374(1), ZN => gl_rom_n_539);
  gl_rom_g35882 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_188(0), B1 => gl_rom_n_20, B2 => gl_rom_rom_186(0), ZN => gl_rom_n_538);
  gl_rom_g35883 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_368(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_371(1), ZN => gl_rom_n_537);
  gl_rom_g35884 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_338(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_343(1), ZN => gl_rom_n_536);
  gl_rom_g35885 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_185(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_189(0), ZN => gl_rom_n_535);
  gl_rom_g35886 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_337(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_341(1), ZN => gl_rom_n_534);
  gl_rom_g35887 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_644(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_646(0), ZN => gl_rom_n_533);
  gl_rom_g35888 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_340(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_339(1), ZN => gl_rom_n_532);
  gl_rom_g35889 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_184(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_187(0), ZN => gl_rom_n_531);
  gl_rom_g35890 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_336(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_342(1), ZN => gl_rom_n_530);
  gl_rom_g35891 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_600(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_601(0), ZN => gl_rom_n_529);
  gl_rom_g35892 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_378(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_383(1), ZN => gl_rom_n_528);
  gl_rom_g35893 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_642(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_647(0), ZN => gl_rom_n_527);
  gl_rom_g35894 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_380(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_382(1), ZN => gl_rom_n_526);
  gl_rom_g35895 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_169(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_173(0), ZN => gl_rom_n_525);
  gl_rom_g35896 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_172(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_174(0), ZN => gl_rom_n_524);
  gl_rom_g35897 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_381(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_379(1), ZN => gl_rom_n_523);
  gl_rom_g35898 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_376(1), B1 => gl_rom_n_21, B2 => gl_rom_rom_377(1), ZN => gl_rom_n_522);
  gl_rom_g35899 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_362(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_367(1), ZN => gl_rom_n_521);
  gl_rom_g35900 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_640(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_643(0), ZN => gl_rom_n_520);
  gl_rom_g35901 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_170(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_171(0), ZN => gl_rom_n_519);
  gl_rom_g35902 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_364(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_366(1), ZN => gl_rom_n_518);
  gl_rom_g35903 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_168(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_175(0), ZN => gl_rom_n_517);
  gl_rom_g35904 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_365(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_363(1), ZN => gl_rom_n_516);
  gl_rom_g35905 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_360(1), B1 => gl_rom_n_21, B2 => gl_rom_rom_361(1), ZN => gl_rom_n_515);
  gl_rom_g35906 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_922(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_927(0), ZN => gl_rom_n_514);
  gl_rom_g35907 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_334(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_335(1), ZN => gl_rom_n_513);
  gl_rom_g35908 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_332(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_330(1), ZN => gl_rom_n_512);
  gl_rom_g35909 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_154(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_159(0), ZN => gl_rom_n_511);
  gl_rom_g35910 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_610(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_615(0), ZN => gl_rom_n_510);
  gl_rom_g35911 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_329(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_333(1), ZN => gl_rom_n_509);
  gl_rom_g35912 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_328(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_331(1), ZN => gl_rom_n_508);
  gl_rom_g35913 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_156(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_158(0), ZN => gl_rom_n_507);
  gl_rom_g35914 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_326(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_327(1), ZN => gl_rom_n_506);
  gl_rom_g35915 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_561(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_565(0), ZN => gl_rom_n_505);
  gl_rom_g35916 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_157(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_155(0), ZN => gl_rom_n_504);
  gl_rom_g35917 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_324(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_322(1), ZN => gl_rom_n_503);
  gl_rom_g35918 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_564(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_566(0), ZN => gl_rom_n_502);
  gl_rom_g35919 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_152(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_153(0), ZN => gl_rom_n_501);
  gl_rom_g35920 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_321(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_325(1), ZN => gl_rom_n_500);
  gl_rom_g35921 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_320(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_323(1), ZN => gl_rom_n_499);
  gl_rom_g35922 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_609(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_613(0), ZN => gl_rom_n_498);
  gl_rom_g35923 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_122(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_127(1), ZN => gl_rom_n_497);
  gl_rom_g35924 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_166(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_167(0), ZN => gl_rom_n_496);
  gl_rom_g35925 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_121(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_125(1), ZN => gl_rom_n_495);
  gl_rom_g35926 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_124(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_126(1), ZN => gl_rom_n_494);
  gl_rom_g35927 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_562(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_563(0), ZN => gl_rom_n_493);
  gl_rom_g35928 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_164(0), B1 => gl_rom_n_20, B2 => gl_rom_rom_162(0), ZN => gl_rom_n_492);
  gl_rom_g35929 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_120(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_123(1), ZN => gl_rom_n_491);
  gl_rom_g35930 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_920(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_923(0), ZN => gl_rom_n_490);
  gl_rom_g35931 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_110(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_111(1), ZN => gl_rom_n_489);
  gl_rom_g35932 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_161(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_165(0), ZN => gl_rom_n_488);
  gl_rom_g35933 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_560(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_567(0), ZN => gl_rom_n_487);
  gl_rom_g35934 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_108(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_106(1), ZN => gl_rom_n_486);
  gl_rom_g35935 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_160(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_163(0), ZN => gl_rom_n_485);
  gl_rom_g35936 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_105(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_109(1), ZN => gl_rom_n_484);
  gl_rom_g35937 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_104(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_107(1), ZN => gl_rom_n_483);
  gl_rom_g35938 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_1002(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_1003(0), ZN => gl_rom_n_482);
  gl_rom_g35939 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_94(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_95(1), ZN => gl_rom_n_481);
  gl_rom_g35940 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_612(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_611(0), ZN => gl_rom_n_480);
  gl_rom_g35941 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_92(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_90(1), ZN => gl_rom_n_479);
  gl_rom_g35942 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_178(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_183(0), ZN => gl_rom_n_478);
  gl_rom_g35943 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_89(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_93(1), ZN => gl_rom_n_477);
  gl_rom_g35944 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_608(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_614(0), ZN => gl_rom_n_476);
  gl_rom_g35945 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_180(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_182(0), ZN => gl_rom_n_475);
  gl_rom_g35946 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_88(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_91(1), ZN => gl_rom_n_474);
  gl_rom_g35947 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_529(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_533(0), ZN => gl_rom_n_473);
  gl_rom_g35948 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_97(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_101(1), ZN => gl_rom_n_472);
  gl_rom_g35949 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_532(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_534(0), ZN => gl_rom_n_471);
  gl_rom_g35950 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_100(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_102(1), ZN => gl_rom_n_470);
  gl_rom_g35951 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_181(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_179(0), ZN => gl_rom_n_469);
  gl_rom_g35952 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_98(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_99(1), ZN => gl_rom_n_468);
  gl_rom_g35953 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_176(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_177(0), ZN => gl_rom_n_467);
  gl_rom_g35954 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_96(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_103(1), ZN => gl_rom_n_466);
  gl_rom_g35955 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_114(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_119(1), ZN => gl_rom_n_465);
  gl_rom_g35956 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_146(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_151(0), ZN => gl_rom_n_464);
  gl_rom_g35957 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_113(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_117(1), ZN => gl_rom_n_463);
  gl_rom_g35958 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_530(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_535(0), ZN => gl_rom_n_462);
  gl_rom_g35959 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_116(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_115(1), ZN => gl_rom_n_461);
  gl_rom_g35960 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_148(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_150(0), ZN => gl_rom_n_460);
  gl_rom_g35961 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_112(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_118(1), ZN => gl_rom_n_459);
  gl_rom_g35962 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_82(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_87(1), ZN => gl_rom_n_458);
  gl_rom_g35963 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_149(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_147(0), ZN => gl_rom_n_457);
  gl_rom_g35964 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_84(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_86(1), ZN => gl_rom_n_456);
  gl_rom_g35965 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_1000(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_1007(0), ZN => gl_rom_n_455);
  gl_rom_g35966 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_528(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_531(0), ZN => gl_rom_n_454);
  gl_rom_g35967 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_85(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_83(1), ZN => gl_rom_n_453);
  gl_rom_g35968 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_144(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_145(0), ZN => gl_rom_n_452);
  gl_rom_g35969 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_80(1), B1 => gl_rom_n_21, B2 => gl_rom_rom_81(1), ZN => gl_rom_n_451);
  gl_rom_g35970 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_930(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_935(0), ZN => gl_rom_n_450);
  gl_rom_g35971 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_73(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_77(1), ZN => gl_rom_n_449);
  gl_rom_g35972 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_138(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_143(0), ZN => gl_rom_n_448);
  gl_rom_g35973 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_76(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_78(1), ZN => gl_rom_n_447);
  gl_rom_g35974 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_74(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_75(1), ZN => gl_rom_n_446);
  gl_rom_g35975 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_625(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_629(0), ZN => gl_rom_n_445);
  gl_rom_g35976 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_140(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_142(0), ZN => gl_rom_n_444);
  gl_rom_g35977 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_72(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_79(1), ZN => gl_rom_n_443);
  gl_rom_g35978 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_538(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_543(0), ZN => gl_rom_n_442);
  gl_rom_g35979 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_70(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_71(1), ZN => gl_rom_n_441);
  gl_rom_g35980 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_141(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_139(0), ZN => gl_rom_n_440);
  gl_rom_g35981 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_68(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_66(1), ZN => gl_rom_n_439);
  gl_rom_g35982 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_136(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_137(0), ZN => gl_rom_n_438);
  gl_rom_g35983 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_65(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_69(1), ZN => gl_rom_n_437);
  gl_rom_g35984 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_64(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_67(1), ZN => gl_rom_n_436);
  gl_rom_g35985 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_537(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_541(0), ZN => gl_rom_n_435);
  gl_rom_g35986 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_130(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_135(0), ZN => gl_rom_n_434);
  gl_rom_g35987 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_182(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_183(1), ZN => gl_rom_n_433);
  gl_rom_g35988 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_628(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_630(0), ZN => gl_rom_n_432);
  gl_rom_g35989 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_180(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_178(1), ZN => gl_rom_n_431);
  gl_rom_g35990 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_129(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_133(0), ZN => gl_rom_n_430);
  gl_rom_g35991 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_177(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_181(1), ZN => gl_rom_n_429);
  gl_rom_g35992 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_540(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_539(0), ZN => gl_rom_n_428);
  gl_rom_g35993 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_176(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_179(1), ZN => gl_rom_n_427);
  gl_rom_g35994 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_132(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_134(0), ZN => gl_rom_n_426);
  gl_rom_g35995 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_986(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_991(0), ZN => gl_rom_n_425);
  gl_rom_g35996 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_536(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_542(0), ZN => gl_rom_n_424);
  gl_rom_g35997 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_150(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_151(1), ZN => gl_rom_n_423);
  gl_rom_g35998 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_148(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_146(1), ZN => gl_rom_n_422);
  gl_rom_g35999 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_128(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_131(0), ZN => gl_rom_n_421);
  gl_rom_g36000 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_145(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_149(1), ZN => gl_rom_n_420);
  gl_rom_g36001 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_929(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_933(0), ZN => gl_rom_n_419);
  gl_rom_g36002 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_144(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_147(1), ZN => gl_rom_n_418);
  gl_rom_g36003 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_158(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_159(1), ZN => gl_rom_n_417);
  gl_rom_g36004 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_626(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_627(0), ZN => gl_rom_n_416);
  gl_rom_g36005 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_156(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_154(1), ZN => gl_rom_n_415);
  gl_rom_g36006 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_58(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_63(0), ZN => gl_rom_n_414);
  gl_rom_g36007 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_153(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_157(1), ZN => gl_rom_n_413);
  gl_rom_g36008 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_545(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_549(0), ZN => gl_rom_n_412);
  gl_rom_g36009 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_152(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_155(1), ZN => gl_rom_n_411);
  gl_rom_g36010 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_57(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_61(0), ZN => gl_rom_n_410);
  gl_rom_g36011 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_162(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_167(1), ZN => gl_rom_n_409);
  gl_rom_g36012 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_164(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_166(1), ZN => gl_rom_n_408);
  gl_rom_g36013 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_60(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_62(0), ZN => gl_rom_n_407);
  gl_rom_g36014 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_56(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_59(0), ZN => gl_rom_n_406);
  gl_rom_g36015 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_165(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_163(1), ZN => gl_rom_n_405);
  gl_rom_g36016 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_160(1), B1 => gl_rom_n_21, B2 => gl_rom_rom_161(1), ZN => gl_rom_n_404);
  gl_rom_g36017 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_548(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_550(0), ZN => gl_rom_n_403);
  gl_rom_g36018 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_190(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_191(1), ZN => gl_rom_n_402);
  gl_rom_g36019 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_624(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_631(0), ZN => gl_rom_n_401);
  gl_rom_g36020 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_46(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_47(0), ZN => gl_rom_n_400);
  gl_rom_g36021 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_188(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_186(1), ZN => gl_rom_n_399);
  gl_rom_g36022 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_546(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_551(0), ZN => gl_rom_n_398);
  gl_rom_g36023 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_185(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_189(1), ZN => gl_rom_n_397);
  gl_rom_g36024 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_44(0), B1 => gl_rom_n_20, B2 => gl_rom_rom_42(0), ZN => gl_rom_n_396);
  gl_rom_g36025 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_184(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_187(1), ZN => gl_rom_n_395);
  gl_rom_g36026 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_170(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_175(1), ZN => gl_rom_n_394);
  gl_rom_g36027 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_544(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_547(0), ZN => gl_rom_n_393);
  gl_rom_g36028 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_41(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_45(0), ZN => gl_rom_n_392);
  gl_rom_g36029 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_172(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_174(1), ZN => gl_rom_n_391);
  gl_rom_g36030 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_40(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_43(0), ZN => gl_rom_n_390);
  gl_rom_g36031 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_173(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_171(1), ZN => gl_rom_n_389);
  gl_rom_g36032 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_168(1), B1 => gl_rom_n_21, B2 => gl_rom_rom_169(1), ZN => gl_rom_n_388);
  gl_rom_g36033 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_1013(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_1011(0), ZN => gl_rom_n_387);
  gl_rom_g36034 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_932(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_931(0), ZN => gl_rom_n_386);
  gl_rom_g36035 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_142(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_143(1), ZN => gl_rom_n_385);
  gl_rom_g36036 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_594(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_599(0), ZN => gl_rom_n_384);
  gl_rom_g36037 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_140(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_138(1), ZN => gl_rom_n_383);
  gl_rom_g36038 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_50(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_55(0), ZN => gl_rom_n_382);
  gl_rom_g36039 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_137(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_141(1), ZN => gl_rom_n_381);
  gl_rom_g36040 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_52(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_54(0), ZN => gl_rom_n_380);
  gl_rom_g36041 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_136(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_139(1), ZN => gl_rom_n_379);
  gl_rom_g36042 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_570(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_575(0), ZN => gl_rom_n_378);
  gl_rom_g36043 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_134(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_135(1), ZN => gl_rom_n_377);
  gl_rom_g36044 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_53(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_51(0), ZN => gl_rom_n_376);
  gl_rom_g36045 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_132(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_130(1), ZN => gl_rom_n_375);
  gl_rom_g36046 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_572(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_574(0), ZN => gl_rom_n_374);
  gl_rom_g36047 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_48(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_49(0), ZN => gl_rom_n_373);
  gl_rom_g36048 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_129(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_133(1), ZN => gl_rom_n_372);
  gl_rom_g36049 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_128(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_131(1), ZN => gl_rom_n_371);
  gl_rom_g36050 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_593(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_597(0), ZN => gl_rom_n_370);
  gl_rom_g36051 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_62(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_63(1), ZN => gl_rom_n_369);
  gl_rom_g36052 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_17(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_21(0), ZN => gl_rom_n_368);
  gl_rom_g36053 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_60(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_58(1), ZN => gl_rom_n_367);
  gl_rom_g36054 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_57(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_61(1), ZN => gl_rom_n_366);
  gl_rom_g36055 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_20(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_22(0), ZN => gl_rom_n_365);
  gl_rom_g36056 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_56(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_59(1), ZN => gl_rom_n_364);
  gl_rom_g36057 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_928(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_934(0), ZN => gl_rom_n_363);
  gl_rom_g36058 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_573(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_571(0), ZN => gl_rom_n_362);
  gl_rom_g36059 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_18(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_19(0), ZN => gl_rom_n_361);
  gl_rom_g36060 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_46(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_47(1), ZN => gl_rom_n_360);
  gl_rom_g36061 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_568(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_569(0), ZN => gl_rom_n_359);
  gl_rom_g36062 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_44(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_42(1), ZN => gl_rom_n_358);
  gl_rom_g36063 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_16(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_23(0), ZN => gl_rom_n_357);
  gl_rom_g36064 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_41(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_45(1), ZN => gl_rom_n_356);
  gl_rom_g36065 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_40(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_43(1), ZN => gl_rom_n_355);
  gl_rom_g36066 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_54(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_55(1), ZN => gl_rom_n_354);
  gl_rom_g36067 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_596(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_598(0), ZN => gl_rom_n_353);
  gl_rom_g36068 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_26(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_31(0), ZN => gl_rom_n_352);
  gl_rom_g36069 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_52(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_50(1), ZN => gl_rom_n_351);
  gl_rom_g36070 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_553(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_557(0), ZN => gl_rom_n_350);
  gl_rom_g36071 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_49(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_53(1), ZN => gl_rom_n_349);
  gl_rom_g36072 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_25(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_29(0), ZN => gl_rom_n_348);
  gl_rom_g36073 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_48(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_51(1), ZN => gl_rom_n_347);
  gl_rom_g36074 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_17(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_21(1), ZN => gl_rom_n_346);
  gl_rom_g36075 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_969(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_973(0), ZN => gl_rom_n_345);
  gl_rom_g36076 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_20(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_22(1), ZN => gl_rom_n_344);
  gl_rom_g36077 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_28(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_27(0), ZN => gl_rom_n_343);
  gl_rom_g36078 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_592(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_595(0), ZN => gl_rom_n_342);
  gl_rom_g36079 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_556(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_558(0), ZN => gl_rom_n_341);
  gl_rom_g36080 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_18(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_19(1), ZN => gl_rom_n_340);
  gl_rom_g36081 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_24(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_30(0), ZN => gl_rom_n_339);
  gl_rom_g36082 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_16(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_23(1), ZN => gl_rom_n_338);
  gl_rom_g36083 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_30(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_31(1), ZN => gl_rom_n_337);
  gl_rom_g36084 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_34(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_39(0), ZN => gl_rom_n_336);
  gl_rom_g36085 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_28(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_26(1), ZN => gl_rom_n_335);
  gl_rom_g36086 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_36(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_38(0), ZN => gl_rom_n_334);
  gl_rom_g36087 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_25(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_29(1), ZN => gl_rom_n_333);
  gl_rom_g36088 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_24(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_27(1), ZN => gl_rom_n_332);
  gl_rom_g36089 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_554(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_555(0), ZN => gl_rom_n_331);
  gl_rom_g36090 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_34(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_39(1), ZN => gl_rom_n_330);
  gl_rom_g36091 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_552(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_559(0), ZN => gl_rom_n_329);
  gl_rom_g36092 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_37(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_35(0), ZN => gl_rom_n_328);
  gl_rom_g36093 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_33(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_37(1), ZN => gl_rom_n_327);
  gl_rom_g36094 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_988(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_990(0), ZN => gl_rom_n_326);
  gl_rom_g36095 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_32(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_33(0), ZN => gl_rom_n_325);
  gl_rom_g36096 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_36(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_38(1), ZN => gl_rom_n_324);
  gl_rom_g36097 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_32(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_35(1), ZN => gl_rom_n_323);
  gl_rom_g36098 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_910(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_911(0), ZN => gl_rom_n_322);
  gl_rom_g36099 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_9(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_13(1), ZN => gl_rom_n_321);
  gl_rom_g36100 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_14(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_15(0), ZN => gl_rom_n_320);
  gl_rom_g36101 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_12(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_14(1), ZN => gl_rom_n_319);
  gl_rom_g36102 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_10(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_11(1), ZN => gl_rom_n_318);
  gl_rom_g36103 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_586(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_591(0), ZN => gl_rom_n_317);
  gl_rom_g36104 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_12(0), B1 => gl_rom_n_20, B2 => gl_rom_rom_10(0), ZN => gl_rom_n_316);
  gl_rom_g36105 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_8(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_15(1), ZN => gl_rom_n_315);
  gl_rom_g36106 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_526(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_527(0), ZN => gl_rom_n_314);
  gl_rom_g36107 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_524(0), B1 => gl_rom_n_20, B2 => gl_rom_rom_522(0), ZN => gl_rom_n_313);
  gl_rom_g36108 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_9(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_13(0), ZN => gl_rom_n_312);
  gl_rom_g36109 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_2(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_7(1), ZN => gl_rom_n_311);
  gl_rom_g36110 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_1(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_5(1), ZN => gl_rom_n_310);
  gl_rom_g36111 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_588(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_590(0), ZN => gl_rom_n_309);
  gl_rom_g36112 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_8(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_11(0), ZN => gl_rom_n_308);
  gl_rom_g36113 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_4(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_6(1), ZN => gl_rom_n_307);
  gl_rom_g36114 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_0(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_3(1), ZN => gl_rom_n_306);
  gl_rom_g36115 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_1(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_5(0), ZN => gl_rom_n_305);
  gl_rom_g36116 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_521(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_525(0), ZN => gl_rom_n_304);
  gl_rom_g36117 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_4(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_6(0), ZN => gl_rom_n_303);
  gl_rom_g36118 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_908(0), B1 => gl_rom_n_20, B2 => gl_rom_rom_906(0), ZN => gl_rom_n_302);
  gl_rom_g36119 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_520(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_523(0), ZN => gl_rom_n_301);
  gl_rom_g36120 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_2(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_3(0), ZN => gl_rom_n_300);
  gl_rom_g36121 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_0(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_7(0), ZN => gl_rom_n_299);
  gl_rom_g36122 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_589(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_587(0), ZN => gl_rom_n_298);
  gl_rom_g36123 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_513(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_517(0), ZN => gl_rom_n_297);
  gl_rom_g36124 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_516(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_518(0), ZN => gl_rom_n_296);
  gl_rom_g36125 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_894(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_895(1), ZN => gl_rom_n_295);
  gl_rom_g36126 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_353(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_357(1), ZN => gl_rom_n_294);
  gl_rom_g36127 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_584(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_585(0), ZN => gl_rom_n_293);
  gl_rom_g36128 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_889(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_893(1), ZN => gl_rom_n_292);
  gl_rom_g36129 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_514(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_515(0), ZN => gl_rom_n_291);
  gl_rom_g36130 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_888(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_891(1), ZN => gl_rom_n_290);
  gl_rom_g36131 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_972(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_974(0), ZN => gl_rom_n_289);
  gl_rom_g36132 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_905(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_909(0), ZN => gl_rom_n_288);
  gl_rom_g36133 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_878(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_879(1), ZN => gl_rom_n_287);
  gl_rom_g36134 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_512(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_519(0), ZN => gl_rom_n_286);
  gl_rom_g36135 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_876(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_874(1), ZN => gl_rom_n_285);
  gl_rom_g36136 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_873(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_877(1), ZN => gl_rom_n_284);
  gl_rom_g36137 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_872(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_875(1), ZN => gl_rom_n_283);
  gl_rom_g36138 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_578(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_583(0), ZN => gl_rom_n_282);
  gl_rom_g36139 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_580(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_582(0), ZN => gl_rom_n_281);
  gl_rom_g36140 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_862(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_863(1), ZN => gl_rom_n_280);
  gl_rom_g36141 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_904(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_907(0), ZN => gl_rom_n_279);
  gl_rom_g36142 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_860(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_858(1), ZN => gl_rom_n_278);
  gl_rom_g36143 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_506(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_511(0), ZN => gl_rom_n_277);
  gl_rom_g36144 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_857(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_861(1), ZN => gl_rom_n_276);
  gl_rom_g36145 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_505(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_509(0), ZN => gl_rom_n_275);
  gl_rom_g36146 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_856(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_859(1), ZN => gl_rom_n_274);
  gl_rom_g36147 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_870(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_871(1), ZN => gl_rom_n_273);
  gl_rom_g36148 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_868(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_866(1), ZN => gl_rom_n_272);
  gl_rom_g36149 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_989(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_987(0), ZN => gl_rom_n_271);
  gl_rom_g36150 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_581(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_579(0), ZN => gl_rom_n_270);
  gl_rom_g36151 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_508(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_510(0), ZN => gl_rom_n_269);
  gl_rom_g36152 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_865(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_869(1), ZN => gl_rom_n_268);
  gl_rom_g36153 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_864(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_867(1), ZN => gl_rom_n_267);
  gl_rom_g36154 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_504(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_507(0), ZN => gl_rom_n_266);
  gl_rom_g36155 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_970(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_971(0), ZN => gl_rom_n_265);
  gl_rom_g36156 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_886(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_887(1), ZN => gl_rom_n_264);
  gl_rom_g36157 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_884(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_882(1), ZN => gl_rom_n_263);
  gl_rom_g36158 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_576(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_577(0), ZN => gl_rom_n_262);
  gl_rom_g36159 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_494(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_495(0), ZN => gl_rom_n_261);
  gl_rom_g36160 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_881(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_885(1), ZN => gl_rom_n_260);
  gl_rom_g36161 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_492(0), B1 => gl_rom_n_20, B2 => gl_rom_rom_490(0), ZN => gl_rom_n_259);
  gl_rom_g36162 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_880(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_883(1), ZN => gl_rom_n_258);
  gl_rom_g36163 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_968(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_975(0), ZN => gl_rom_n_257);
  gl_rom_g36164 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_854(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_855(1), ZN => gl_rom_n_256);
  gl_rom_g36165 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_852(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_850(1), ZN => gl_rom_n_255);
  gl_rom_g36166 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_489(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_493(0), ZN => gl_rom_n_254);
  gl_rom_g36167 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_897(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_901(0), ZN => gl_rom_n_253);
  gl_rom_g36168 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_849(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_853(1), ZN => gl_rom_n_252);
  gl_rom_g36169 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_848(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_851(1), ZN => gl_rom_n_251);
  gl_rom_g36170 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_488(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_491(0), ZN => gl_rom_n_250);
  gl_rom_g36171 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_900(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_902(0), ZN => gl_rom_n_249);
  gl_rom_g36172 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_841(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_845(1), ZN => gl_rom_n_248);
  gl_rom_g36173 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_844(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_846(1), ZN => gl_rom_n_247);
  gl_rom_g36174 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_478(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_479(0), ZN => gl_rom_n_246);
  gl_rom_g36175 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_842(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_843(1), ZN => gl_rom_n_245);
  gl_rom_g36176 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_754(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_759(0), ZN => gl_rom_n_244);
  gl_rom_g36177 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_840(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_847(1), ZN => gl_rom_n_243);
  gl_rom_g36178 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_476(0), B1 => gl_rom_n_20, B2 => gl_rom_rom_474(0), ZN => gl_rom_n_242);
  gl_rom_g36179 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_833(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_837(1), ZN => gl_rom_n_241);
  gl_rom_g36180 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_836(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_838(1), ZN => gl_rom_n_240);
  gl_rom_g36181 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_473(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_477(0), ZN => gl_rom_n_239);
  gl_rom_g36182 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_834(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_835(1), ZN => gl_rom_n_238);
  gl_rom_g36183 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_472(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_475(0), ZN => gl_rom_n_237);
  gl_rom_g36184 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_832(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_839(1), ZN => gl_rom_n_236);
  gl_rom_g36185 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_753(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_757(0), ZN => gl_rom_n_235);
  gl_rom_g36186 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_601(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_605(1), ZN => gl_rom_n_234);
  gl_rom_g36187 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_604(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_606(1), ZN => gl_rom_n_233);
  gl_rom_g36188 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_482(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_487(0), ZN => gl_rom_n_232);
  gl_rom_g36189 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_756(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_755(0), ZN => gl_rom_n_231);
  gl_rom_g36190 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_602(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_603(1), ZN => gl_rom_n_230);
  gl_rom_g36191 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_600(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_607(1), ZN => gl_rom_n_229);
  gl_rom_g36192 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_481(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_485(0), ZN => gl_rom_n_228);
  gl_rom_g36193 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_752(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_758(0), ZN => gl_rom_n_227);
  gl_rom_g36194 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_609(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_613(1), ZN => gl_rom_n_226);
  gl_rom_g36195 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_484(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_486(0), ZN => gl_rom_n_225);
  gl_rom_g36196 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_612(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_614(1), ZN => gl_rom_n_224);
  gl_rom_g36197 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_898(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_899(0), ZN => gl_rom_n_223);
  gl_rom_g36198 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_480(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_483(0), ZN => gl_rom_n_222);
  gl_rom_g36199 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_610(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_611(1), ZN => gl_rom_n_221);
  gl_rom_g36200 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_608(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_615(1), ZN => gl_rom_n_220);
  gl_rom_g36201 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_626(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_631(1), ZN => gl_rom_n_219);
  gl_rom_g36202 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_896(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_903(0), ZN => gl_rom_n_218);
  gl_rom_g36203 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_625(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_629(1), ZN => gl_rom_n_217);
  gl_rom_g36204 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_722(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_727(0), ZN => gl_rom_n_216);
  gl_rom_g36205 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_502(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_503(0), ZN => gl_rom_n_215);
  gl_rom_g36206 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_628(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_630(1), ZN => gl_rom_n_214);
  gl_rom_g36207 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_624(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_627(1), ZN => gl_rom_n_213);
  gl_rom_g36208 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_500(0), B1 => gl_rom_n_20, B2 => gl_rom_rom_498(0), ZN => gl_rom_n_212);
  gl_rom_g36209 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_724(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_726(0), ZN => gl_rom_n_211);
  gl_rom_g36210 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_593(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_597(1), ZN => gl_rom_n_210);
  gl_rom_g36211 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_596(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_598(1), ZN => gl_rom_n_209);
  gl_rom_g36212 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_497(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_501(0), ZN => gl_rom_n_208);
  gl_rom_g36213 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_594(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_599(1), ZN => gl_rom_n_207);
  gl_rom_g36214 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_592(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_595(1), ZN => gl_rom_n_206);
  gl_rom_g36215 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_496(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_499(0), ZN => gl_rom_n_205);
  gl_rom_g36216 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_634(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_639(1), ZN => gl_rom_n_204);
  gl_rom_g36217 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_984(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_985(0), ZN => gl_rom_n_203);
  gl_rom_g36218 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_1008(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_1009(0), ZN => gl_rom_n_202);
  gl_rom_g36219 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_465(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_469(0), ZN => gl_rom_n_201);
  gl_rom_g36220 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_636(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_638(1), ZN => gl_rom_n_200);
  gl_rom_g36221 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_725(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_723(0), ZN => gl_rom_n_199);
  gl_rom_g36222 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_637(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_635(1), ZN => gl_rom_n_198);
  gl_rom_g36223 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_468(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_470(0), ZN => gl_rom_n_197);
  gl_rom_g36224 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_632(1), B1 => gl_rom_n_21, B2 => gl_rom_rom_633(1), ZN => gl_rom_n_196);
  gl_rom_g36225 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_962(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_967(0), ZN => gl_rom_n_195);
  gl_rom_g36226 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_618(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_623(1), ZN => gl_rom_n_194);
  gl_rom_g36227 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_720(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_721(0), ZN => gl_rom_n_193);
  gl_rom_g36228 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_617(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_621(1), ZN => gl_rom_n_192);
  gl_rom_g36229 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_466(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_467(0), ZN => gl_rom_n_191);
  gl_rom_g36230 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_620(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_619(1), ZN => gl_rom_n_190);
  gl_rom_g36231 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_464(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_471(0), ZN => gl_rom_n_189);
  gl_rom_g36232 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_616(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_622(1), ZN => gl_rom_n_188);
  gl_rom_g36233 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_590(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_591(1), ZN => gl_rom_n_187);
  gl_rom_g36234 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_588(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_586(1), ZN => gl_rom_n_186);
  gl_rom_g36235 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_462(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_463(0), ZN => gl_rom_n_185);
  gl_rom_g36236 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_585(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_589(1), ZN => gl_rom_n_184);
  gl_rom_g36237 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_730(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_735(0), ZN => gl_rom_n_183);
  gl_rom_g36238 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_460(0), B1 => gl_rom_n_20, B2 => gl_rom_rom_458(0), ZN => gl_rom_n_182);
  gl_rom_g36239 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_584(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_587(1), ZN => gl_rom_n_181);
  gl_rom_g36240 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_964(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_966(0), ZN => gl_rom_n_180);
  gl_rom_g36241 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_577(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_581(1), ZN => gl_rom_n_179);
  gl_rom_g36242 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_729(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_733(0), ZN => gl_rom_n_178);
  gl_rom_g36243 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_580(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_582(1), ZN => gl_rom_n_177);
  gl_rom_g36244 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_457(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_461(0), ZN => gl_rom_n_176);
  gl_rom_g36245 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_857(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_861(0), ZN => gl_rom_n_175);
  gl_rom_g36246 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_578(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_579(1), ZN => gl_rom_n_174);
  gl_rom_g36247 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_576(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_583(1), ZN => gl_rom_n_173);
  gl_rom_g36248 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_456(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_459(0), ZN => gl_rom_n_172);
  gl_rom_g36249 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_860(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_862(0), ZN => gl_rom_n_171);
  gl_rom_g36250 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_761(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_765(1), ZN => gl_rom_n_170);
  gl_rom_g36251 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_732(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_731(0), ZN => gl_rom_n_169);
  gl_rom_g36252 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_454(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_455(0), ZN => gl_rom_n_168);
  gl_rom_g36253 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_764(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_766(1), ZN => gl_rom_n_167);
  gl_rom_g36254 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_452(0), B1 => gl_rom_n_20, B2 => gl_rom_rom_450(0), ZN => gl_rom_n_166);
  gl_rom_g36255 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_762(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_767(1), ZN => gl_rom_n_165);
  gl_rom_g36256 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_760(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_763(1), ZN => gl_rom_n_164);
  gl_rom_g36257 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_728(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_734(0), ZN => gl_rom_n_163);
  gl_rom_g36258 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_449(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_453(0), ZN => gl_rom_n_162);
  gl_rom_g36259 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_746(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_751(1), ZN => gl_rom_n_161);
  gl_rom_g36260 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_748(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_750(1), ZN => gl_rom_n_160);
  gl_rom_g36261 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_448(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_451(0), ZN => gl_rom_n_159);
  gl_rom_g36262 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_749(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_747(1), ZN => gl_rom_n_158);
  gl_rom_g36263 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_744(1), B1 => gl_rom_n_21, B2 => gl_rom_rom_745(1), ZN => gl_rom_n_157);
  gl_rom_g36264 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_753(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_757(1), ZN => gl_rom_n_156);
  gl_rom_g36265 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_756(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_758(1), ZN => gl_rom_n_155);
  gl_rom_g36266 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_738(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_743(0), ZN => gl_rom_n_154);
  gl_rom_g36267 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_446(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_447(0), ZN => gl_rom_n_153);
  gl_rom_g36268 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_754(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_759(1), ZN => gl_rom_n_152);
  gl_rom_g36269 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_858(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_859(0), ZN => gl_rom_n_151);
  gl_rom_g36270 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_752(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_755(1), ZN => gl_rom_n_150);
  gl_rom_g36271 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_444(0), B1 => gl_rom_n_20, B2 => gl_rom_rom_442(0), ZN => gl_rom_n_149);
  gl_rom_g36272 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_740(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_742(0), ZN => gl_rom_n_148);
  gl_rom_g36273 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_721(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_725(1), ZN => gl_rom_n_147);
  gl_rom_g36274 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_724(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_726(1), ZN => gl_rom_n_146);
  gl_rom_g36275 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_441(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_445(0), ZN => gl_rom_n_145);
  gl_rom_g36276 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_965(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_963(0), ZN => gl_rom_n_144);
  gl_rom_g36277 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_722(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_723(1), ZN => gl_rom_n_143);
  gl_rom_g36278 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_720(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_727(1), ZN => gl_rom_n_142);
  gl_rom_g36279 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_440(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_443(0), ZN => gl_rom_n_141);
  gl_rom_g36280 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_856(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_863(0), ZN => gl_rom_n_140);
  gl_rom_g36281 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_741(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_739(0), ZN => gl_rom_n_139);
  gl_rom_g36282 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_730(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_735(1), ZN => gl_rom_n_138);
  gl_rom_g36283 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_732(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_734(1), ZN => gl_rom_n_137);
  gl_rom_g36284 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_425(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_429(0), ZN => gl_rom_n_136);
  gl_rom_g36285 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_733(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_731(1), ZN => gl_rom_n_135);
  gl_rom_g36286 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_428(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_430(0), ZN => gl_rom_n_134);
  gl_rom_g36287 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_728(1), B1 => gl_rom_n_21, B2 => gl_rom_rom_729(1), ZN => gl_rom_n_133);
  gl_rom_g36288 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_736(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_737(0), ZN => gl_rom_n_132);
  gl_rom_g36289 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_738(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_743(1), ZN => gl_rom_n_131);
  gl_rom_g36290 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_426(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_427(0), ZN => gl_rom_n_130);
  gl_rom_g36291 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_740(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_742(1), ZN => gl_rom_n_129);
  gl_rom_g36292 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_741(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_739(1), ZN => gl_rom_n_128);
  gl_rom_g36293 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_424(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_431(0), ZN => gl_rom_n_127);
  gl_rom_g36294 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_736(1), B1 => gl_rom_n_21, B2 => gl_rom_rom_737(1), ZN => gl_rom_n_126);
  gl_rom_g36295 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_714(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_719(1), ZN => gl_rom_n_125);
  gl_rom_g36296 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_716(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_718(1), ZN => gl_rom_n_124);
  gl_rom_g36297 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_414(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_415(0), ZN => gl_rom_n_123);
  gl_rom_g36298 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_761(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_765(0), ZN => gl_rom_n_122);
  gl_rom_g36299 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_717(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_715(1), ZN => gl_rom_n_121);
  gl_rom_g36300 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_712(1), B1 => gl_rom_n_21, B2 => gl_rom_rom_713(1), ZN => gl_rom_n_120);
  gl_rom_g36301 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_865(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_869(0), ZN => gl_rom_n_119);
  gl_rom_g36302 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_412(0), B1 => gl_rom_n_20, B2 => gl_rom_rom_410(0), ZN => gl_rom_n_118);
  gl_rom_g36303 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_706(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_711(1), ZN => gl_rom_n_117);
  gl_rom_g36304 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_960(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_961(0), ZN => gl_rom_n_116);
  gl_rom_g36305 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_705(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_709(1), ZN => gl_rom_n_115);
  gl_rom_g36306 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_764(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_766(0), ZN => gl_rom_n_114);
  gl_rom_g36307 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_409(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_413(0), ZN => gl_rom_n_113);
  gl_rom_g36308 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_408(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_411(0), ZN => gl_rom_n_112);
  gl_rom_g36309 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_708(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_707(1), ZN => gl_rom_n_111);
  gl_rom_g36310 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_704(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_710(1), ZN => gl_rom_n_110);
  gl_rom_g36311 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_868(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_870(0), ZN => gl_rom_n_109);
  gl_rom_g36312 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_826(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_831(1), ZN => gl_rom_n_108);
  gl_rom_g36313 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_762(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_763(0), ZN => gl_rom_n_107);
  gl_rom_g36314 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_422(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_423(0), ZN => gl_rom_n_106);
  gl_rom_g36315 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_825(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_829(1), ZN => gl_rom_n_105);
  gl_rom_g36316 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_420(0), B1 => gl_rom_n_20, B2 => gl_rom_rom_418(0), ZN => gl_rom_n_104);
  gl_rom_g36317 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_828(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_830(1), ZN => gl_rom_n_103);
  gl_rom_g36318 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_824(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_827(1), ZN => gl_rom_n_102);
  gl_rom_g36319 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_760(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_767(0), ZN => gl_rom_n_101);
  gl_rom_g36320 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_809(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_813(1), ZN => gl_rom_n_100);
  gl_rom_g36321 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_417(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_421(0), ZN => gl_rom_n_99);
  gl_rom_g36322 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_812(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_814(1), ZN => gl_rom_n_98);
  gl_rom_g36323 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_416(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_419(0), ZN => gl_rom_n_97);
  gl_rom_g36324 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_810(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_815(1), ZN => gl_rom_n_96);
  gl_rom_g36325 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_808(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_811(1), ZN => gl_rom_n_95);
  gl_rom_g36326 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_798(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_799(1), ZN => gl_rom_n_94);
  gl_rom_g36327 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_994(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_999(0), ZN => gl_rom_n_93);
  gl_rom_g36328 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_796(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_794(1), ZN => gl_rom_n_92);
  gl_rom_g36329 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_866(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_867(0), ZN => gl_rom_n_91);
  gl_rom_g36330 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_438(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_439(0), ZN => gl_rom_n_90);
  gl_rom_g36331 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_746(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_751(0), ZN => gl_rom_n_89);
  gl_rom_g36332 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_793(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_797(1), ZN => gl_rom_n_88);
  gl_rom_g36333 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_792(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_795(1), ZN => gl_rom_n_87);
  gl_rom_g36334 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_436(0), B1 => gl_rom_n_20, B2 => gl_rom_rom_434(0), ZN => gl_rom_n_86);
  gl_rom_g36335 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_748(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_750(0), ZN => gl_rom_n_85);
  gl_rom_g36336 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_806(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_807(1), ZN => gl_rom_n_84);
  gl_rom_g36337 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_804(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_802(1), ZN => gl_rom_n_83);
  gl_rom_g36338 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_433(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_437(0), ZN => gl_rom_n_82);
  gl_rom_g36339 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_801(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_805(1), ZN => gl_rom_n_81);
  gl_rom_g36340 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_800(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_803(1), ZN => gl_rom_n_80);
  gl_rom_g36341 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_432(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_435(0), ZN => gl_rom_n_79);
  gl_rom_g36342 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_1010(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_1015(0), ZN => gl_rom_n_78);
  gl_rom_g36343 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_749(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_747(0), ZN => gl_rom_n_77);
  gl_rom_g36344 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_818(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_823(1), ZN => gl_rom_n_76);
  gl_rom_g36345 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_864(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_871(0), ZN => gl_rom_n_75);
  gl_rom_g36346 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_406(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_407(0), ZN => gl_rom_n_74);
  gl_rom_g36347 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_817(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_821(1), ZN => gl_rom_n_73);
  gl_rom_g36348 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_996(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_998(0), ZN => gl_rom_n_72);
  gl_rom_g36349 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_820(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_822(1), ZN => gl_rom_n_71);
  gl_rom_g36350 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_404(0), B1 => gl_rom_n_20, B2 => gl_rom_rom_402(0), ZN => gl_rom_n_70);
  gl_rom_g36351 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_816(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_819(1), ZN => gl_rom_n_69);
  gl_rom_g36352 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_744(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_745(0), ZN => gl_rom_n_68);
  gl_rom_g36353 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_790(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_791(1), ZN => gl_rom_n_67);
  gl_rom_g36354 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_788(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_786(1), ZN => gl_rom_n_66);
  gl_rom_g36355 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_401(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_405(0), ZN => gl_rom_n_65);
  gl_rom_g36356 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_785(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_789(1), ZN => gl_rom_n_64);
  gl_rom_g36357 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_400(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_403(0), ZN => gl_rom_n_63);
  gl_rom_g36358 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_784(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_787(1), ZN => gl_rom_n_62);
  gl_rom_g36359 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_777(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_781(1), ZN => gl_rom_n_61);
  gl_rom_g36360 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_780(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_782(1), ZN => gl_rom_n_60);
  gl_rom_g36361 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_398(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_399(0), ZN => gl_rom_n_59);
  gl_rom_g36362 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_714(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_719(0), ZN => gl_rom_n_58);
  gl_rom_g36363 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_778(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_779(1), ZN => gl_rom_n_57);
  gl_rom_g36364 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_396(0), B1 => gl_rom_n_20, B2 => gl_rom_rom_394(0), ZN => gl_rom_n_56);
  gl_rom_g36365 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_776(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_783(1), ZN => gl_rom_n_55);
  gl_rom_g36366 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_774(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_775(1), ZN => gl_rom_n_54);
  gl_rom_g36367 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_716(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_718(0), ZN => gl_rom_n_53);
  gl_rom_g36368 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_393(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_397(0), ZN => gl_rom_n_52);
  gl_rom_g36369 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_772(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_770(1), ZN => gl_rom_n_51);
  gl_rom_g36370 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_881(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_885(0), ZN => gl_rom_n_50);
  gl_rom_g36371 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_392(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_395(0), ZN => gl_rom_n_49);
  gl_rom_g36372 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_769(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_773(1), ZN => gl_rom_n_48);
  gl_rom_g36373 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_768(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_771(1), ZN => gl_rom_n_47);
  gl_rom_g36374 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_954(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_959(0), ZN => gl_rom_n_46);
  gl_rom_g36375 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_884(0), B1 => gl_rom_n_16, B2 => gl_rom_rom_886(0), ZN => gl_rom_n_45);
  gl_rom_g36376 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_717(0), B1 => gl_rom_n_15, B2 => gl_rom_rom_715(0), ZN => gl_rom_n_44);
  gl_rom_g36377 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_1014(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_1015(1), ZN => gl_rom_n_43);
  gl_rom_g36378 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_390(0), B1 => gl_rom_n_17, B2 => gl_rom_rom_391(0), ZN => gl_rom_n_42);
  gl_rom_g36379 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_1012(1), B1 => gl_rom_n_20, B2 => gl_rom_rom_1010(1), ZN => gl_rom_n_41);
  gl_rom_g36380 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_388(0), B1 => gl_rom_n_20, B2 => gl_rom_rom_386(0), ZN => gl_rom_n_40);
  gl_rom_g36381 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_1009(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_1013(1), ZN => gl_rom_n_39);
  gl_rom_g36382 : AN2D1BWP7T port map(A1 => gl_rom_n_13, A2 => gl_sig_e(8), Z => gl_rom_n_38);
  gl_rom_g36383 : INR2D1BWP7T port map(A1 => gl_sig_e(8), B1 => gl_rom_n_1, ZN => gl_rom_n_37);
  gl_rom_g36384 : INR2D1BWP7T port map(A1 => gl_sig_e(8), B1 => gl_rom_n_2, ZN => gl_rom_n_36);
  gl_rom_g36385 : NR2D1BWP7T port map(A1 => gl_rom_n_1, A2 => gl_sig_e(8), ZN => gl_rom_n_35);
  gl_rom_g36386 : NR2D1BWP7T port map(A1 => gl_rom_n_9, A2 => gl_sig_e(8), ZN => gl_rom_n_34);
  gl_rom_g36387 : NR2D1BWP7T port map(A1 => gl_rom_n_2, A2 => gl_sig_e(8), ZN => gl_rom_n_33);
  gl_rom_g36388 : INR2D1BWP7T port map(A1 => gl_rom_n_13, B1 => gl_sig_e(8), ZN => gl_rom_n_32);
  gl_rom_g36389 : INR2D1BWP7T port map(A1 => gl_sig_e(8), B1 => gl_rom_n_9, ZN => gl_rom_n_31);
  gl_rom_g36390 : AN2D1BWP7T port map(A1 => gl_rom_n_8, A2 => gl_sig_e(4), Z => gl_rom_n_30);
  gl_rom_g36391 : NR2D1BWP7T port map(A1 => gl_rom_n_7, A2 => gl_sig_e(4), ZN => gl_rom_n_29);
  gl_rom_g36392 : AN2D1BWP7T port map(A1 => gl_rom_n_4, A2 => gl_sig_e(4), Z => gl_rom_n_28);
  gl_rom_g36393 : INR2D1BWP7T port map(A1 => gl_sig_e(4), B1 => gl_rom_n_11, ZN => gl_rom_n_27);
  gl_rom_g36394 : NR2D1BWP7T port map(A1 => gl_rom_n_11, A2 => gl_sig_e(4), ZN => gl_rom_n_26);
  gl_rom_g36395 : AN2D1BWP7T port map(A1 => gl_rom_n_14, A2 => gl_sig_e(4), Z => gl_rom_n_25);
  gl_rom_g36396 : INR2D1BWP7T port map(A1 => gl_rom_n_14, B1 => gl_sig_e(4), ZN => gl_rom_n_24);
  gl_rom_g36397 : NR2D1BWP7T port map(A1 => gl_rom_n_5, A2 => gl_sig_e(4), ZN => gl_rom_n_23);
  gl_rom_g36398 : AN2D4BWP7T port map(A1 => gl_rom_n_3, A2 => gl_sig_e(2), Z => gl_rom_n_22);
  gl_rom_g36399 : AN2D4BWP7T port map(A1 => gl_rom_n_3, A2 => gl_rom_n_0, Z => gl_rom_n_21);
  gl_rom_g36400 : AN2D4BWP7T port map(A1 => gl_rom_n_10, A2 => gl_rom_n_0, Z => gl_rom_n_20);
  gl_rom_g36401 : AN2D4BWP7T port map(A1 => gl_rom_n_6, A2 => gl_rom_n_0, Z => gl_rom_n_19);
  gl_rom_g36402 : AN2D4BWP7T port map(A1 => gl_rom_n_6, A2 => gl_sig_e(2), Z => gl_rom_n_18);
  gl_rom_g36403 : AN2D4BWP7T port map(A1 => gl_rom_n_12, A2 => gl_sig_e(2), Z => gl_rom_n_17);
  gl_rom_g36404 : AN2D4BWP7T port map(A1 => gl_rom_n_10, A2 => gl_sig_e(2), Z => gl_rom_n_16);
  gl_rom_g36405 : AN2D4BWP7T port map(A1 => gl_rom_n_12, A2 => gl_rom_n_0, Z => gl_rom_n_15);
  gl_rom_g36406 : NR2XD0BWP7T port map(A1 => gl_sig_e(5), A2 => gl_sig_e(3), ZN => gl_rom_n_14);
  gl_rom_g36407 : NR2D0BWP7T port map(A1 => gl_sig_e(7), A2 => gl_sig_e(6), ZN => gl_rom_n_13);
  gl_rom_g36408 : AN2D1BWP7T port map(A1 => gl_sig_e(1), A2 => gl_sig_e(0), Z => gl_rom_n_12);
  gl_rom_g36409 : ND2D1BWP7T port map(A1 => gl_sig_e(3), A2 => gl_sig_e(5), ZN => gl_rom_n_11);
  gl_rom_g36410 : INR2D1BWP7T port map(A1 => gl_sig_e(1), B1 => gl_sig_e(0), ZN => gl_rom_n_10);
  gl_rom_g36411 : CKND2D1BWP7T port map(A1 => gl_sig_e(7), A2 => gl_sig_e(6), ZN => gl_rom_n_9);
  gl_rom_g36412 : INVD0BWP7T port map(I => gl_rom_n_7, ZN => gl_rom_n_8);
  gl_rom_g36413 : INVD0BWP7T port map(I => gl_rom_n_4, ZN => gl_rom_n_5);
  gl_rom_g36414 : IND2D1BWP7T port map(A1 => gl_sig_e(5), B1 => gl_sig_e(3), ZN => gl_rom_n_7);
  gl_rom_g36415 : NR2D1BWP7T port map(A1 => gl_sig_e(1), A2 => gl_sig_e(0), ZN => gl_rom_n_6);
  gl_rom_g36416 : INR2D1BWP7T port map(A1 => gl_sig_e(5), B1 => gl_sig_e(3), ZN => gl_rom_n_4);
  gl_rom_g36417 : INR2D1BWP7T port map(A1 => gl_sig_e(0), B1 => gl_sig_e(1), ZN => gl_rom_n_3);
  gl_rom_g36418 : IND2D1BWP7T port map(A1 => gl_sig_e(7), B1 => gl_sig_e(6), ZN => gl_rom_n_2);
  gl_rom_g36419 : IND2D1BWP7T port map(A1 => gl_sig_e(6), B1 => gl_sig_e(7), ZN => gl_rom_n_1);
  gl_rom_g36420 : INVD2BWP7T port map(I => gl_sig_e(2), ZN => gl_rom_n_0);
  gl_ram_g13798 : MOAI22D0BWP7T port map(A1 => gl_ram_n_1059, A2 => gl_ram_n_1027, B1 => gl_ram_n_1055, B2 => gl_ram_n_1027, ZN => gl_sig_ram(2));
  gl_ram_g13799 : MOAI22D0BWP7T port map(A1 => gl_ram_n_1058, A2 => gl_ram_n_1027, B1 => gl_ram_n_1054, B2 => gl_ram_n_1027, ZN => gl_sig_ram(0));
  gl_ram_g13800 : MOAI22D0BWP7T port map(A1 => gl_ram_n_1057, A2 => gl_ram_n_1027, B1 => gl_ram_n_1056, B2 => gl_ram_n_1027, ZN => gl_sig_ram(1));
  gl_ram_g13801 : AN4D0BWP7T port map(A1 => gl_ram_n_1052, A2 => gl_ram_n_1053, A3 => gl_ram_n_1033, A4 => gl_ram_n_1043, Z => gl_ram_n_1059);
  gl_ram_g13802 : AN4D0BWP7T port map(A1 => gl_ram_n_1051, A2 => gl_ram_n_1050, A3 => gl_ram_n_1032, A4 => gl_ram_n_1040, Z => gl_ram_n_1058);
  gl_ram_g13803 : AN4D0BWP7T port map(A1 => gl_ram_n_1048, A2 => gl_ram_n_1049, A3 => gl_ram_n_1031, A4 => gl_ram_n_1037, Z => gl_ram_n_1057);
  gl_ram_g13804 : ND4D0BWP7T port map(A1 => gl_ram_n_1035, A2 => gl_ram_n_1042, A3 => gl_ram_n_1039, A4 => gl_ram_n_1044, ZN => gl_ram_n_1056);
  gl_ram_g13805 : ND4D0BWP7T port map(A1 => gl_ram_n_1034, A2 => gl_ram_n_1041, A3 => gl_ram_n_1045, A4 => gl_ram_n_1047, ZN => gl_ram_n_1055);
  gl_ram_g13806 : ND4D0BWP7T port map(A1 => gl_ram_n_1038, A2 => gl_ram_n_1036, A3 => gl_ram_n_1046, A4 => gl_ram_n_1030, ZN => gl_ram_n_1054);
  gl_ram_g13807 : AOI22D0BWP7T port map(A1 => gl_ram_n_1028, A2 => gl_ram_ram_96(2), B1 => gl_ram_n_803, B2 => gl_ram_ram_97(2), ZN => gl_ram_n_1053);
  gl_ram_g13808 : AOI22D0BWP7T port map(A1 => gl_ram_n_1029, A2 => gl_ram_ram_98(2), B1 => gl_ram_n_802, B2 => gl_ram_ram_99(2), ZN => gl_ram_n_1052);
  gl_ram_g13809 : AOI22D0BWP7T port map(A1 => gl_ram_n_1029, A2 => gl_ram_ram_98(0), B1 => gl_ram_n_802, B2 => gl_ram_ram_99(0), ZN => gl_ram_n_1051);
  gl_ram_g13810 : AOI22D0BWP7T port map(A1 => gl_ram_n_1028, A2 => gl_ram_ram_96(0), B1 => gl_ram_n_803, B2 => gl_ram_ram_97(0), ZN => gl_ram_n_1050);
  gl_ram_g13811 : AOI22D0BWP7T port map(A1 => gl_ram_n_1028, A2 => gl_ram_ram_96(1), B1 => gl_ram_n_803, B2 => gl_ram_ram_97(1), ZN => gl_ram_n_1049);
  gl_ram_g13812 : AOI22D0BWP7T port map(A1 => gl_ram_n_1029, A2 => gl_ram_ram_98(1), B1 => gl_ram_n_802, B2 => gl_ram_ram_99(1), ZN => gl_ram_n_1048);
  gl_ram_g13813 : AOI22D0BWP7T port map(A1 => gl_ram_n_1020, A2 => gl_ram_n_982, B1 => gl_ram_n_1026, B2 => gl_ram_n_989, ZN => gl_ram_n_1047);
  gl_ram_g13814 : AOI22D0BWP7T port map(A1 => gl_ram_n_1022, A2 => gl_ram_n_990, B1 => gl_ram_n_1021, B2 => gl_ram_n_983, ZN => gl_ram_n_1046);
  gl_ram_g13815 : AOI22D0BWP7T port map(A1 => gl_ram_n_1022, A2 => gl_ram_n_1006, B1 => gl_ram_n_1021, B2 => gl_ram_n_974, ZN => gl_ram_n_1045);
  gl_ram_g13816 : AOI22D0BWP7T port map(A1 => gl_ram_n_1020, A2 => gl_ram_n_1007, B1 => gl_ram_n_1026, B2 => gl_ram_n_999, ZN => gl_ram_n_1044);
  gl_ram_g13817 : AOI22D0BWP7T port map(A1 => gl_ram_n_1025, A2 => gl_ram_n_997, B1 => gl_ram_n_1024, B2 => gl_ram_n_1004, ZN => gl_ram_n_1043);
  gl_ram_g13818 : AOI22D0BWP7T port map(A1 => gl_ram_n_1025, A2 => gl_ram_n_996, B1 => gl_ram_n_1018, B2 => gl_ram_n_998, ZN => gl_ram_n_1042);
  gl_ram_g13819 : AOI22D0BWP7T port map(A1 => gl_ram_n_1025, A2 => gl_ram_n_992, B1 => gl_ram_n_1018, B2 => gl_ram_n_994, ZN => gl_ram_n_1041);
  gl_ram_g13820 : AOI22D0BWP7T port map(A1 => gl_ram_n_1025, A2 => gl_ram_n_988, B1 => gl_ram_n_1024, B2 => gl_ram_n_981, ZN => gl_ram_n_1040);
  gl_ram_g13821 : AOI22D0BWP7T port map(A1 => gl_ram_n_1022, A2 => gl_ram_n_1000, B1 => gl_ram_n_1021, B2 => gl_ram_n_1001, ZN => gl_ram_n_1039);
  gl_ram_g13822 : AOI22D0BWP7T port map(A1 => gl_ram_n_1019, A2 => gl_ram_n_977, B1 => gl_ram_n_1024, B2 => gl_ram_n_979, ZN => gl_ram_n_1038);
  gl_ram_g13823 : AOI22D0BWP7T port map(A1 => gl_ram_n_1025, A2 => gl_ram_n_976, B1 => gl_ram_n_1024, B2 => gl_ram_n_980, ZN => gl_ram_n_1037);
  gl_ram_g13824 : AOI22D0BWP7T port map(A1 => gl_ram_n_1025, A2 => gl_ram_n_973, B1 => gl_ram_n_1018, B2 => gl_ram_n_975, ZN => gl_ram_n_1036);
  gl_ram_g13825 : AOI22D0BWP7T port map(A1 => gl_ram_n_1019, A2 => gl_ram_n_1003, B1 => gl_ram_n_1024, B2 => gl_ram_n_1005, ZN => gl_ram_n_1035);
  gl_ram_g13826 : AOI22D0BWP7T port map(A1 => gl_ram_n_1019, A2 => gl_ram_n_1008, B1 => gl_ram_n_1024, B2 => gl_ram_n_1002, ZN => gl_ram_n_1034);
  gl_ram_g13827 : AOI22D0BWP7T port map(A1 => gl_ram_n_1019, A2 => gl_ram_n_978, B1 => gl_ram_n_1018, B2 => gl_ram_n_995, ZN => gl_ram_n_1033);
  gl_ram_g13828 : AOI22D0BWP7T port map(A1 => gl_ram_n_1019, A2 => gl_ram_n_991, B1 => gl_ram_n_1018, B2 => gl_ram_n_993, ZN => gl_ram_n_1032);
  gl_ram_g13829 : AOI22D0BWP7T port map(A1 => gl_ram_n_1019, A2 => gl_ram_n_984, B1 => gl_ram_n_1018, B2 => gl_ram_n_987, ZN => gl_ram_n_1031);
  gl_ram_g13830 : AOI22D0BWP7T port map(A1 => gl_ram_n_1020, A2 => gl_ram_n_985, B1 => gl_ram_n_1026, B2 => gl_ram_n_986, ZN => gl_ram_n_1030);
  gl_ram_g13831 : NR2D0BWP7T port map(A1 => gl_ram_n_1023, A2 => gl_ram_n_824, ZN => gl_ram_n_1029);
  gl_ram_g13832 : NR2D0BWP7T port map(A1 => gl_ram_n_1023, A2 => gl_ram_n_822, ZN => gl_ram_n_1028);
  gl_ram_g13835 : XNR2D1BWP7T port map(A1 => gl_ram_n_1015, A2 => gl_sig_y(3), ZN => gl_ram_n_1027);
  gl_ram_g13836 : INVD0BWP7T port map(I => gl_ram_n_1023, ZN => gl_ram_n_1022);
  gl_ram_g13837 : NR2D0BWP7T port map(A1 => gl_ram_n_1016, A2 => gl_ram_n_1013, ZN => gl_ram_n_1026);
  gl_ram_g13838 : INR2D0BWP7T port map(A1 => gl_ram_n_1012, B1 => gl_ram_n_1017, ZN => gl_ram_n_1025);
  gl_ram_g13839 : NR2D0BWP7T port map(A1 => gl_ram_n_1017, A2 => gl_ram_n_1013, ZN => gl_ram_n_1024);
  gl_ram_g13840 : ND2D0BWP7T port map(A1 => gl_ram_n_1017, A2 => gl_ram_n_1012, ZN => gl_ram_n_1023);
  gl_ram_g13841 : NR2D0BWP7T port map(A1 => gl_ram_n_1016, A2 => gl_ram_n_1014, ZN => gl_ram_n_1021);
  gl_ram_g13842 : NR2D0BWP7T port map(A1 => gl_ram_n_1016, A2 => gl_ram_n_1011, ZN => gl_ram_n_1020);
  gl_ram_g13843 : NR2D0BWP7T port map(A1 => gl_ram_n_1017, A2 => gl_ram_n_1014, ZN => gl_ram_n_1019);
  gl_ram_g13844 : NR2D0BWP7T port map(A1 => gl_ram_n_1017, A2 => gl_ram_n_1011, ZN => gl_ram_n_1018);
  gl_ram_g13845 : CKND1BWP7T port map(I => gl_ram_n_1017, ZN => gl_ram_n_1016);
  gl_ram_g13846 : FA1D0BWP7T port map(A => gl_ram_n_806, B => gl_sig_y(2), CI => gl_ram_n_1009, CO => gl_ram_n_1015, S => gl_ram_n_1017);
  gl_ram_g13847 : IND2D0BWP7T port map(A1 => gl_ram_n_1010, B1 => gl_ram_n_972, ZN => gl_ram_n_1014);
  gl_ram_g13848 : ND2D0BWP7T port map(A1 => gl_ram_n_1010, A2 => gl_ram_n_972, ZN => gl_ram_n_1013);
  gl_ram_g13849 : NR2D0BWP7T port map(A1 => gl_ram_n_1010, A2 => gl_ram_n_972, ZN => gl_ram_n_1012);
  gl_ram_g13850 : IND2D0BWP7T port map(A1 => gl_ram_n_972, B1 => gl_ram_n_1010, ZN => gl_ram_n_1011);
  gl_ram_g13851 : FA1D0BWP7T port map(A => gl_ram_n_807, B => gl_ram_n_808, CI => gl_ram_n_971, CO => gl_ram_n_1009, S => gl_ram_n_1010);
  gl_ram_g13852 : ND4D0BWP7T port map(A1 => gl_ram_n_925, A2 => gl_ram_n_917, A3 => gl_ram_n_927, A4 => gl_ram_n_922, ZN => gl_ram_n_1008);
  gl_ram_g13853 : ND4D0BWP7T port map(A1 => gl_ram_n_959, A2 => gl_ram_n_956, A3 => gl_ram_n_960, A4 => gl_ram_n_958, ZN => gl_ram_n_1007);
  gl_ram_g13854 : ND4D0BWP7T port map(A1 => gl_ram_n_955, A2 => gl_ram_n_948, A3 => gl_ram_n_957, A4 => gl_ram_n_952, ZN => gl_ram_n_1006);
  gl_ram_g13855 : ND4D0BWP7T port map(A1 => gl_ram_n_953, A2 => gl_ram_n_949, A3 => gl_ram_n_954, A4 => gl_ram_n_951, ZN => gl_ram_n_1005);
  gl_ram_g13856 : ND4D0BWP7T port map(A1 => gl_ram_n_943, A2 => gl_ram_n_930, A3 => gl_ram_n_950, A4 => gl_ram_n_937, ZN => gl_ram_n_1004);
  gl_ram_g13857 : ND4D0BWP7T port map(A1 => gl_ram_n_944, A2 => gl_ram_n_941, A3 => gl_ram_n_947, A4 => gl_ram_n_946, ZN => gl_ram_n_1003);
  gl_ram_g13858 : ND4D0BWP7T port map(A1 => gl_ram_n_936, A2 => gl_ram_n_932, A3 => gl_ram_n_942, A4 => gl_ram_n_940, ZN => gl_ram_n_1002);
  gl_ram_g13859 : ND4D0BWP7T port map(A1 => gl_ram_n_935, A2 => gl_ram_n_934, A3 => gl_ram_n_939, A4 => gl_ram_n_938, ZN => gl_ram_n_1001);
  gl_ram_g13860 : ND4D0BWP7T port map(A1 => gl_ram_n_929, A2 => gl_ram_n_926, A3 => gl_ram_n_931, A4 => gl_ram_n_928, ZN => gl_ram_n_1000);
  gl_ram_g13861 : ND4D0BWP7T port map(A1 => gl_ram_n_964, A2 => gl_ram_n_962, A3 => gl_ram_n_967, A4 => gl_ram_n_966, ZN => gl_ram_n_999);
  gl_ram_g13862 : ND4D0BWP7T port map(A1 => gl_ram_n_923, A2 => gl_ram_n_919, A3 => gl_ram_n_924, A4 => gl_ram_n_921, ZN => gl_ram_n_998);
  gl_ram_g13863 : ND4D0BWP7T port map(A1 => gl_ram_n_908, A2 => gl_ram_n_901, A3 => gl_ram_n_918, A4 => gl_ram_n_906, ZN => gl_ram_n_997);
  gl_ram_g13864 : ND4D0BWP7T port map(A1 => gl_ram_n_914, A2 => gl_ram_n_910, A3 => gl_ram_n_915, A4 => gl_ram_n_913, ZN => gl_ram_n_996);
  gl_ram_g13865 : ND4D0BWP7T port map(A1 => gl_ram_n_970, A2 => gl_ram_n_865, A3 => gl_ram_n_909, A4 => gl_ram_n_884, ZN => gl_ram_n_995);
  gl_ram_g13866 : ND4D0BWP7T port map(A1 => gl_ram_n_907, A2 => gl_ram_n_904, A3 => gl_ram_n_912, A4 => gl_ram_n_911, ZN => gl_ram_n_994);
  gl_ram_g13867 : ND4D0BWP7T port map(A1 => gl_ram_n_902, A2 => gl_ram_n_900, A3 => gl_ram_n_905, A4 => gl_ram_n_903, ZN => gl_ram_n_993);
  gl_ram_g13868 : ND4D0BWP7T port map(A1 => gl_ram_n_895, A2 => gl_ram_n_890, A3 => gl_ram_n_827, A4 => gl_ram_n_892, ZN => gl_ram_n_992);
  gl_ram_g13869 : ND4D0BWP7T port map(A1 => gl_ram_n_896, A2 => gl_ram_n_893, A3 => gl_ram_n_897, A4 => gl_ram_n_894, ZN => gl_ram_n_991);
  gl_ram_g13870 : ND4D0BWP7T port map(A1 => gl_ram_n_854, A2 => gl_ram_n_852, A3 => gl_ram_n_856, A4 => gl_ram_n_853, ZN => gl_ram_n_990);
  gl_ram_g13871 : ND4D0BWP7T port map(A1 => gl_ram_n_880, A2 => gl_ram_n_868, A3 => gl_ram_n_886, A4 => gl_ram_n_876, ZN => gl_ram_n_989);
  gl_ram_g13872 : ND4D0BWP7T port map(A1 => gl_ram_n_883, A2 => gl_ram_n_881, A3 => gl_ram_n_885, A4 => gl_ram_n_882, ZN => gl_ram_n_988);
  gl_ram_g13873 : ND4D0BWP7T port map(A1 => gl_ram_n_875, A2 => gl_ram_n_869, A3 => gl_ram_n_878, A4 => gl_ram_n_872, ZN => gl_ram_n_987);
  gl_ram_g13874 : ND4D0BWP7T port map(A1 => gl_ram_n_874, A2 => gl_ram_n_873, A3 => gl_ram_n_879, A4 => gl_ram_n_877, ZN => gl_ram_n_986);
  gl_ram_g13875 : ND4D0BWP7T port map(A1 => gl_ram_n_870, A2 => gl_ram_n_866, A3 => gl_ram_n_871, A4 => gl_ram_n_867, ZN => gl_ram_n_985);
  gl_ram_g13876 : ND4D0BWP7T port map(A1 => gl_ram_n_861, A2 => gl_ram_n_855, A3 => gl_ram_n_863, A4 => gl_ram_n_857, ZN => gl_ram_n_984);
  gl_ram_g13877 : ND4D0BWP7T port map(A1 => gl_ram_n_862, A2 => gl_ram_n_859, A3 => gl_ram_n_864, A4 => gl_ram_n_860, ZN => gl_ram_n_983);
  gl_ram_g13878 : ND4D0BWP7T port map(A1 => gl_ram_n_851, A2 => gl_ram_n_920, A3 => gl_ram_n_858, A4 => gl_ram_n_845, ZN => gl_ram_n_982);
  gl_ram_g13879 : ND4D0BWP7T port map(A1 => gl_ram_n_889, A2 => gl_ram_n_887, A3 => gl_ram_n_891, A4 => gl_ram_n_888, ZN => gl_ram_n_981);
  gl_ram_g13880 : ND4D0BWP7T port map(A1 => gl_ram_n_847, A2 => gl_ram_n_842, A3 => gl_ram_n_850, A4 => gl_ram_n_933, ZN => gl_ram_n_980);
  gl_ram_g13881 : ND4D0BWP7T port map(A1 => gl_ram_n_916, A2 => gl_ram_n_846, A3 => gl_ram_n_849, A4 => gl_ram_n_848, ZN => gl_ram_n_979);
  gl_ram_g13882 : ND4D0BWP7T port map(A1 => gl_ram_n_899, A2 => gl_ram_n_961, A3 => gl_ram_n_968, A4 => gl_ram_n_836, ZN => gl_ram_n_978);
  gl_ram_g13883 : ND4D0BWP7T port map(A1 => gl_ram_n_843, A2 => gl_ram_n_840, A3 => gl_ram_n_844, A4 => gl_ram_n_841, ZN => gl_ram_n_977);
  gl_ram_g13884 : ND4D0BWP7T port map(A1 => gl_ram_n_945, A2 => gl_ram_n_898, A3 => gl_ram_n_839, A4 => gl_ram_n_835, ZN => gl_ram_n_976);
  gl_ram_g13885 : ND4D0BWP7T port map(A1 => gl_ram_n_834, A2 => gl_ram_n_833, A3 => gl_ram_n_838, A4 => gl_ram_n_837, ZN => gl_ram_n_975);
  gl_ram_g13886 : ND4D0BWP7T port map(A1 => gl_ram_n_969, A2 => gl_ram_n_963, A3 => gl_ram_n_831, A4 => gl_ram_n_965, ZN => gl_ram_n_974);
  gl_ram_g13887 : ND4D0BWP7T port map(A1 => gl_ram_n_830, A2 => gl_ram_n_828, A3 => gl_ram_n_832, A4 => gl_ram_n_829, ZN => gl_ram_n_973);
  gl_ram_g13888 : FA1D0BWP7T port map(A => gl_ram_n_809, B => gl_sig_y(2), CI => gl_ram_n_814, CO => gl_ram_n_971, S => gl_ram_n_972);
  gl_ram_g13889 : AOI22D0BWP7T port map(A1 => gl_ram_ram_80(2), A2 => gl_ram_n_823, B1 => gl_ram_ram_83(2), B2 => gl_ram_n_817, ZN => gl_ram_n_970);
  gl_ram_g13890 : AOI22D0BWP7T port map(A1 => gl_ram_ram_41(2), A2 => gl_ram_n_821, B1 => gl_ram_ram_42(2), B2 => gl_ram_n_825, ZN => gl_ram_n_969);
  gl_ram_g13891 : AOI22D0BWP7T port map(A1 => gl_ram_ram_78(2), A2 => gl_ram_n_826, B1 => gl_ram_ram_79(2), B2 => gl_ram_n_820, ZN => gl_ram_n_968);
  gl_ram_g13892 : AOI22D0BWP7T port map(A1 => gl_ram_ram_62(1), A2 => gl_ram_n_826, B1 => gl_ram_ram_63(1), B2 => gl_ram_n_820, ZN => gl_ram_n_967);
  gl_ram_g13893 : AOI22D0BWP7T port map(A1 => gl_ram_ram_60(1), A2 => gl_ram_n_819, B1 => gl_ram_ram_61(1), B2 => gl_ram_n_818, ZN => gl_ram_n_966);
  gl_ram_g13894 : AOI22D0BWP7T port map(A1 => gl_ram_ram_44(2), A2 => gl_ram_n_819, B1 => gl_ram_ram_45(2), B2 => gl_ram_n_818, ZN => gl_ram_n_965);
  gl_ram_g13895 : AOI22D0BWP7T port map(A1 => gl_ram_ram_57(1), A2 => gl_ram_n_821, B1 => gl_ram_ram_58(1), B2 => gl_ram_n_825, ZN => gl_ram_n_964);
  gl_ram_g13896 : AOI22D0BWP7T port map(A1 => gl_ram_ram_40(2), A2 => gl_ram_n_823, B1 => gl_ram_ram_43(2), B2 => gl_ram_n_817, ZN => gl_ram_n_963);
  gl_ram_g13897 : AOI22D0BWP7T port map(A1 => gl_ram_ram_56(1), A2 => gl_ram_n_823, B1 => gl_ram_ram_59(1), B2 => gl_ram_n_817, ZN => gl_ram_n_962);
  gl_ram_g13898 : AOI22D0BWP7T port map(A1 => gl_ram_ram_72(2), A2 => gl_ram_n_823, B1 => gl_ram_ram_75(2), B2 => gl_ram_n_817, ZN => gl_ram_n_961);
  gl_ram_g13899 : AOI22D0BWP7T port map(A1 => gl_ram_ram_54(1), A2 => gl_ram_n_826, B1 => gl_ram_ram_55(1), B2 => gl_ram_n_820, ZN => gl_ram_n_960);
  gl_ram_g13900 : AOI22D0BWP7T port map(A1 => gl_ram_ram_49(1), A2 => gl_ram_n_821, B1 => gl_ram_ram_50(1), B2 => gl_ram_n_825, ZN => gl_ram_n_959);
  gl_ram_g13901 : AOI22D0BWP7T port map(A1 => gl_ram_ram_52(1), A2 => gl_ram_n_819, B1 => gl_ram_ram_53(1), B2 => gl_ram_n_818, ZN => gl_ram_n_958);
  gl_ram_g13902 : AOI22D0BWP7T port map(A1 => gl_ram_ram_38(2), A2 => gl_ram_n_826, B1 => gl_ram_ram_39(2), B2 => gl_ram_n_820, ZN => gl_ram_n_957);
  gl_ram_g13903 : AOI22D0BWP7T port map(A1 => gl_ram_ram_48(1), A2 => gl_ram_n_823, B1 => gl_ram_ram_51(1), B2 => gl_ram_n_817, ZN => gl_ram_n_956);
  gl_ram_g13904 : AOI22D0BWP7T port map(A1 => gl_ram_ram_33(2), A2 => gl_ram_n_821, B1 => gl_ram_ram_34(2), B2 => gl_ram_n_825, ZN => gl_ram_n_955);
  gl_ram_g13905 : AOI22D0BWP7T port map(A1 => gl_ram_ram_30(1), A2 => gl_ram_n_826, B1 => gl_ram_ram_31(1), B2 => gl_ram_n_820, ZN => gl_ram_n_954);
  gl_ram_g13906 : AOI22D0BWP7T port map(A1 => gl_ram_ram_24(1), A2 => gl_ram_n_823, B1 => gl_ram_ram_27(1), B2 => gl_ram_n_817, ZN => gl_ram_n_953);
  gl_ram_g13907 : AOI22D0BWP7T port map(A1 => gl_ram_ram_36(2), A2 => gl_ram_n_819, B1 => gl_ram_ram_37(2), B2 => gl_ram_n_818, ZN => gl_ram_n_952);
  gl_ram_g13908 : AOI22D0BWP7T port map(A1 => gl_ram_ram_28(1), A2 => gl_ram_n_819, B1 => gl_ram_ram_29(1), B2 => gl_ram_n_818, ZN => gl_ram_n_951);
  gl_ram_g13909 : AOI22D0BWP7T port map(A1 => gl_ram_ram_94(2), A2 => gl_ram_n_826, B1 => gl_ram_ram_95(2), B2 => gl_ram_n_820, ZN => gl_ram_n_950);
  gl_ram_g13910 : AOI22D0BWP7T port map(A1 => gl_ram_ram_25(1), A2 => gl_ram_n_821, B1 => gl_ram_ram_26(1), B2 => gl_ram_n_825, ZN => gl_ram_n_949);
  gl_ram_g13911 : AOI22D0BWP7T port map(A1 => gl_ram_ram_32(2), A2 => gl_ram_n_823, B1 => gl_ram_ram_35(2), B2 => gl_ram_n_817, ZN => gl_ram_n_948);
  gl_ram_g13912 : AOI22D0BWP7T port map(A1 => gl_ram_ram_14(1), A2 => gl_ram_n_826, B1 => gl_ram_ram_15(1), B2 => gl_ram_n_820, ZN => gl_ram_n_947);
  gl_ram_g13913 : AOI22D0BWP7T port map(A1 => gl_ram_ram_12(1), A2 => gl_ram_n_819, B1 => gl_ram_ram_13(1), B2 => gl_ram_n_818, ZN => gl_ram_n_946);
  gl_ram_g13914 : AOI22D0BWP7T port map(A1 => gl_ram_ram_66(1), A2 => gl_ram_n_825, B1 => gl_ram_ram_67(1), B2 => gl_ram_n_817, ZN => gl_ram_n_945);
  gl_ram_g13915 : AOI22D0BWP7T port map(A1 => gl_ram_ram_10(1), A2 => gl_ram_n_825, B1 => gl_ram_ram_11(1), B2 => gl_ram_n_817, ZN => gl_ram_n_944);
  gl_ram_g13916 : AOI22D0BWP7T port map(A1 => gl_ram_ram_88(2), A2 => gl_ram_n_823, B1 => gl_ram_ram_91(2), B2 => gl_ram_n_817, ZN => gl_ram_n_943);
  gl_ram_g13917 : AOI22D0BWP7T port map(A1 => gl_ram_ram_30(2), A2 => gl_ram_n_826, B1 => gl_ram_ram_31(2), B2 => gl_ram_n_820, ZN => gl_ram_n_942);
  gl_ram_g13918 : AOI22D0BWP7T port map(A1 => gl_ram_ram_8(1), A2 => gl_ram_n_823, B1 => gl_ram_ram_9(1), B2 => gl_ram_n_821, ZN => gl_ram_n_941);
  gl_ram_g13919 : AOI22D0BWP7T port map(A1 => gl_ram_ram_28(2), A2 => gl_ram_n_819, B1 => gl_ram_ram_29(2), B2 => gl_ram_n_818, ZN => gl_ram_n_940);
  gl_ram_g13920 : AOI22D0BWP7T port map(A1 => gl_ram_ram_46(1), A2 => gl_ram_n_826, B1 => gl_ram_ram_47(1), B2 => gl_ram_n_820, ZN => gl_ram_n_939);
  gl_ram_g13921 : AOI22D0BWP7T port map(A1 => gl_ram_ram_44(1), A2 => gl_ram_n_819, B1 => gl_ram_ram_45(1), B2 => gl_ram_n_818, ZN => gl_ram_n_938);
  gl_ram_g13922 : AOI22D0BWP7T port map(A1 => gl_ram_ram_92(2), A2 => gl_ram_n_819, B1 => gl_ram_ram_93(2), B2 => gl_ram_n_818, ZN => gl_ram_n_937);
  gl_ram_g13923 : AOI22D0BWP7T port map(A1 => gl_ram_ram_25(2), A2 => gl_ram_n_821, B1 => gl_ram_ram_26(2), B2 => gl_ram_n_825, ZN => gl_ram_n_936);
  gl_ram_g13924 : AOI22D0BWP7T port map(A1 => gl_ram_ram_41(1), A2 => gl_ram_n_821, B1 => gl_ram_ram_42(1), B2 => gl_ram_n_825, ZN => gl_ram_n_935);
  gl_ram_g13925 : AOI22D0BWP7T port map(A1 => gl_ram_ram_40(1), A2 => gl_ram_n_823, B1 => gl_ram_ram_43(1), B2 => gl_ram_n_817, ZN => gl_ram_n_934);
  gl_ram_g13926 : AOI22D0BWP7T port map(A1 => gl_ram_ram_92(1), A2 => gl_ram_n_819, B1 => gl_ram_ram_93(1), B2 => gl_ram_n_818, ZN => gl_ram_n_933);
  gl_ram_g13927 : AOI22D0BWP7T port map(A1 => gl_ram_ram_24(2), A2 => gl_ram_n_823, B1 => gl_ram_ram_27(2), B2 => gl_ram_n_817, ZN => gl_ram_n_932);
  gl_ram_g13928 : AOI22D0BWP7T port map(A1 => gl_ram_ram_38(1), A2 => gl_ram_n_826, B1 => gl_ram_ram_39(1), B2 => gl_ram_n_820, ZN => gl_ram_n_931);
  gl_ram_g13929 : AOI22D0BWP7T port map(A1 => gl_ram_ram_89(2), A2 => gl_ram_n_821, B1 => gl_ram_ram_90(2), B2 => gl_ram_n_825, ZN => gl_ram_n_930);
  gl_ram_g13930 : AOI22D0BWP7T port map(A1 => gl_ram_ram_33(1), A2 => gl_ram_n_821, B1 => gl_ram_ram_34(1), B2 => gl_ram_n_825, ZN => gl_ram_n_929);
  gl_ram_g13931 : AOI22D0BWP7T port map(A1 => gl_ram_ram_36(1), A2 => gl_ram_n_819, B1 => gl_ram_ram_37(1), B2 => gl_ram_n_818, ZN => gl_ram_n_928);
  gl_ram_g13932 : AOI22D0BWP7T port map(A1 => gl_ram_ram_14(2), A2 => gl_ram_n_826, B1 => gl_ram_ram_15(2), B2 => gl_ram_n_820, ZN => gl_ram_n_927);
  gl_ram_g13933 : AOI22D0BWP7T port map(A1 => gl_ram_ram_32(1), A2 => gl_ram_n_823, B1 => gl_ram_ram_35(1), B2 => gl_ram_n_817, ZN => gl_ram_n_926);
  gl_ram_g13934 : AOI22D0BWP7T port map(A1 => gl_ram_ram_9(2), A2 => gl_ram_n_821, B1 => gl_ram_ram_10(2), B2 => gl_ram_n_825, ZN => gl_ram_n_925);
  gl_ram_g13935 : AOI22D0BWP7T port map(A1 => gl_ram_ram_22(1), A2 => gl_ram_n_826, B1 => gl_ram_ram_23(1), B2 => gl_ram_n_820, ZN => gl_ram_n_924);
  gl_ram_g13936 : AOI22D0BWP7T port map(A1 => gl_ram_ram_16(1), A2 => gl_ram_n_823, B1 => gl_ram_ram_19(1), B2 => gl_ram_n_817, ZN => gl_ram_n_923);
  gl_ram_g13937 : AOI22D0BWP7T port map(A1 => gl_ram_ram_12(2), A2 => gl_ram_n_819, B1 => gl_ram_ram_13(2), B2 => gl_ram_n_818, ZN => gl_ram_n_922);
  gl_ram_g13938 : AOI22D0BWP7T port map(A1 => gl_ram_ram_20(1), A2 => gl_ram_n_819, B1 => gl_ram_ram_21(1), B2 => gl_ram_n_818, ZN => gl_ram_n_921);
  gl_ram_g13939 : AOI22D0BWP7T port map(A1 => gl_ram_ram_49(2), A2 => gl_ram_n_821, B1 => gl_ram_ram_50(2), B2 => gl_ram_n_825, ZN => gl_ram_n_920);
  gl_ram_g13940 : AOI22D0BWP7T port map(A1 => gl_ram_ram_17(1), A2 => gl_ram_n_821, B1 => gl_ram_ram_18(1), B2 => gl_ram_n_825, ZN => gl_ram_n_919);
  gl_ram_g13941 : AOI22D0BWP7T port map(A1 => gl_ram_ram_70(2), A2 => gl_ram_n_826, B1 => gl_ram_ram_71(2), B2 => gl_ram_n_820, ZN => gl_ram_n_918);
  gl_ram_g13942 : AOI22D0BWP7T port map(A1 => gl_ram_ram_8(2), A2 => gl_ram_n_823, B1 => gl_ram_ram_11(2), B2 => gl_ram_n_817, ZN => gl_ram_n_917);
  gl_ram_g13943 : AOI22D0BWP7T port map(A1 => gl_ram_ram_25(0), A2 => gl_ram_n_821, B1 => gl_ram_ram_26(0), B2 => gl_ram_n_825, ZN => gl_ram_n_916);
  gl_ram_g13944 : AOI22D0BWP7T port map(A1 => gl_ram_ram_6(1), A2 => gl_ram_n_826, B1 => gl_ram_ram_7(1), B2 => gl_ram_n_820, ZN => gl_ram_n_915);
  gl_ram_g13945 : AOI22D0BWP7T port map(A1 => gl_ram_ram_1(1), A2 => gl_ram_n_821, B1 => gl_ram_ram_2(1), B2 => gl_ram_n_825, ZN => gl_ram_n_914);
  gl_ram_g13946 : AOI22D0BWP7T port map(A1 => gl_ram_ram_4(1), A2 => gl_ram_n_819, B1 => gl_ram_ram_5(1), B2 => gl_ram_n_818, ZN => gl_ram_n_913);
  gl_ram_g13947 : AOI22D0BWP7T port map(A1 => gl_ram_ram_22(2), A2 => gl_ram_n_826, B1 => gl_ram_ram_23(2), B2 => gl_ram_n_820, ZN => gl_ram_n_912);
  gl_ram_g13948 : AOI22D0BWP7T port map(A1 => gl_ram_ram_20(2), A2 => gl_ram_n_819, B1 => gl_ram_ram_21(2), B2 => gl_ram_n_818, ZN => gl_ram_n_911);
  gl_ram_g13949 : AOI22D0BWP7T port map(A1 => gl_ram_ram_0(1), A2 => gl_ram_n_823, B1 => gl_ram_ram_3(1), B2 => gl_ram_n_817, ZN => gl_ram_n_910);
  gl_ram_g13950 : AOI22D0BWP7T port map(A1 => gl_ram_ram_86(2), A2 => gl_ram_n_826, B1 => gl_ram_ram_87(2), B2 => gl_ram_n_820, ZN => gl_ram_n_909);
  gl_ram_g13951 : AOI22D0BWP7T port map(A1 => gl_ram_ram_65(2), A2 => gl_ram_n_821, B1 => gl_ram_ram_66(2), B2 => gl_ram_n_825, ZN => gl_ram_n_908);
  gl_ram_g13952 : AOI22D0BWP7T port map(A1 => gl_ram_ram_17(2), A2 => gl_ram_n_821, B1 => gl_ram_ram_18(2), B2 => gl_ram_n_825, ZN => gl_ram_n_907);
  gl_ram_g13953 : AOI22D0BWP7T port map(A1 => gl_ram_ram_68(2), A2 => gl_ram_n_819, B1 => gl_ram_ram_69(2), B2 => gl_ram_n_818, ZN => gl_ram_n_906);
  gl_ram_g13954 : AOI22D0BWP7T port map(A1 => gl_ram_ram_86(0), A2 => gl_ram_n_826, B1 => gl_ram_ram_87(0), B2 => gl_ram_n_820, ZN => gl_ram_n_905);
  gl_ram_g13955 : AOI22D0BWP7T port map(A1 => gl_ram_ram_16(2), A2 => gl_ram_n_823, B1 => gl_ram_ram_19(2), B2 => gl_ram_n_817, ZN => gl_ram_n_904);
  gl_ram_g13956 : AOI22D0BWP7T port map(A1 => gl_ram_ram_84(0), A2 => gl_ram_n_819, B1 => gl_ram_ram_85(0), B2 => gl_ram_n_818, ZN => gl_ram_n_903);
  gl_ram_g13957 : AOI22D0BWP7T port map(A1 => gl_ram_ram_81(0), A2 => gl_ram_n_821, B1 => gl_ram_ram_82(0), B2 => gl_ram_n_825, ZN => gl_ram_n_902);
  gl_ram_g13958 : AOI22D0BWP7T port map(A1 => gl_ram_ram_64(2), A2 => gl_ram_n_823, B1 => gl_ram_ram_67(2), B2 => gl_ram_n_817, ZN => gl_ram_n_901);
  gl_ram_g13959 : AOI22D0BWP7T port map(A1 => gl_ram_ram_80(0), A2 => gl_ram_n_823, B1 => gl_ram_ram_83(0), B2 => gl_ram_n_817, ZN => gl_ram_n_900);
  gl_ram_g13960 : AOI22D0BWP7T port map(A1 => gl_ram_ram_73(2), A2 => gl_ram_n_821, B1 => gl_ram_ram_74(2), B2 => gl_ram_n_825, ZN => gl_ram_n_899);
  gl_ram_g13961 : AOI22D0BWP7T port map(A1 => gl_ram_ram_64(1), A2 => gl_ram_n_823, B1 => gl_ram_ram_65(1), B2 => gl_ram_n_821, ZN => gl_ram_n_898);
  gl_ram_g13962 : AOI22D0BWP7T port map(A1 => gl_ram_ram_78(0), A2 => gl_ram_n_826, B1 => gl_ram_ram_79(0), B2 => gl_ram_n_820, ZN => gl_ram_n_897);
  gl_ram_g13963 : AOI22D0BWP7T port map(A1 => gl_ram_ram_72(0), A2 => gl_ram_n_823, B1 => gl_ram_ram_75(0), B2 => gl_ram_n_817, ZN => gl_ram_n_896);
  gl_ram_g13964 : AOI22D0BWP7T port map(A1 => gl_ram_ram_0(2), A2 => gl_ram_n_823, B1 => gl_ram_ram_3(2), B2 => gl_ram_n_817, ZN => gl_ram_n_895);
  gl_ram_g13965 : AOI22D0BWP7T port map(A1 => gl_ram_ram_76(0), A2 => gl_ram_n_819, B1 => gl_ram_ram_77(0), B2 => gl_ram_n_818, ZN => gl_ram_n_894);
  gl_ram_g13966 : AOI22D0BWP7T port map(A1 => gl_ram_ram_73(0), A2 => gl_ram_n_821, B1 => gl_ram_ram_74(0), B2 => gl_ram_n_825, ZN => gl_ram_n_893);
  gl_ram_g13967 : AOI22D0BWP7T port map(A1 => gl_ram_ram_4(2), A2 => gl_ram_n_819, B1 => gl_ram_ram_5(2), B2 => gl_ram_n_818, ZN => gl_ram_n_892);
  gl_ram_g13968 : AOI22D0BWP7T port map(A1 => gl_ram_ram_94(0), A2 => gl_ram_n_826, B1 => gl_ram_ram_95(0), B2 => gl_ram_n_820, ZN => gl_ram_n_891);
  gl_ram_g13969 : AOI22D0BWP7T port map(A1 => gl_ram_ram_1(2), A2 => gl_ram_n_821, B1 => gl_ram_ram_2(2), B2 => gl_ram_n_825, ZN => gl_ram_n_890);
  gl_ram_g13970 : AOI22D0BWP7T port map(A1 => gl_ram_ram_89(0), A2 => gl_ram_n_821, B1 => gl_ram_ram_90(0), B2 => gl_ram_n_825, ZN => gl_ram_n_889);
  gl_ram_g13971 : AOI22D0BWP7T port map(A1 => gl_ram_ram_92(0), A2 => gl_ram_n_819, B1 => gl_ram_ram_93(0), B2 => gl_ram_n_818, ZN => gl_ram_n_888);
  gl_ram_g13972 : AOI22D0BWP7T port map(A1 => gl_ram_ram_88(0), A2 => gl_ram_n_823, B1 => gl_ram_ram_91(0), B2 => gl_ram_n_817, ZN => gl_ram_n_887);
  gl_ram_g13973 : AOI22D0BWP7T port map(A1 => gl_ram_ram_62(2), A2 => gl_ram_n_826, B1 => gl_ram_ram_63(2), B2 => gl_ram_n_820, ZN => gl_ram_n_886);
  gl_ram_g13974 : AOI22D0BWP7T port map(A1 => gl_ram_ram_70(0), A2 => gl_ram_n_826, B1 => gl_ram_ram_71(0), B2 => gl_ram_n_820, ZN => gl_ram_n_885);
  gl_ram_g13975 : AOI22D0BWP7T port map(A1 => gl_ram_ram_84(2), A2 => gl_ram_n_819, B1 => gl_ram_ram_85(2), B2 => gl_ram_n_818, ZN => gl_ram_n_884);
  gl_ram_g13976 : AOI22D0BWP7T port map(A1 => gl_ram_ram_64(0), A2 => gl_ram_n_823, B1 => gl_ram_ram_67(0), B2 => gl_ram_n_817, ZN => gl_ram_n_883);
  gl_ram_g13977 : AOI22D0BWP7T port map(A1 => gl_ram_ram_68(0), A2 => gl_ram_n_819, B1 => gl_ram_ram_69(0), B2 => gl_ram_n_818, ZN => gl_ram_n_882);
  gl_ram_g13978 : AOI22D0BWP7T port map(A1 => gl_ram_ram_65(0), A2 => gl_ram_n_821, B1 => gl_ram_ram_66(0), B2 => gl_ram_n_825, ZN => gl_ram_n_881);
  gl_ram_g13979 : AOI22D0BWP7T port map(A1 => gl_ram_ram_57(2), A2 => gl_ram_n_821, B1 => gl_ram_ram_58(2), B2 => gl_ram_n_825, ZN => gl_ram_n_880);
  gl_ram_g13980 : AOI22D0BWP7T port map(A1 => gl_ram_ram_62(0), A2 => gl_ram_n_826, B1 => gl_ram_ram_63(0), B2 => gl_ram_n_820, ZN => gl_ram_n_879);
  gl_ram_g13981 : AOI22D0BWP7T port map(A1 => gl_ram_ram_86(1), A2 => gl_ram_n_826, B1 => gl_ram_ram_87(1), B2 => gl_ram_n_820, ZN => gl_ram_n_878);
  gl_ram_g13982 : AOI22D0BWP7T port map(A1 => gl_ram_ram_60(0), A2 => gl_ram_n_819, B1 => gl_ram_ram_61(0), B2 => gl_ram_n_818, ZN => gl_ram_n_877);
  gl_ram_g13983 : AOI22D0BWP7T port map(A1 => gl_ram_ram_60(2), A2 => gl_ram_n_819, B1 => gl_ram_ram_61(2), B2 => gl_ram_n_818, ZN => gl_ram_n_876);
  gl_ram_g13984 : AOI22D0BWP7T port map(A1 => gl_ram_ram_81(1), A2 => gl_ram_n_821, B1 => gl_ram_ram_82(1), B2 => gl_ram_n_825, ZN => gl_ram_n_875);
  gl_ram_g13985 : AOI22D0BWP7T port map(A1 => gl_ram_ram_57(0), A2 => gl_ram_n_821, B1 => gl_ram_ram_58(0), B2 => gl_ram_n_825, ZN => gl_ram_n_874);
  gl_ram_g13986 : AOI22D0BWP7T port map(A1 => gl_ram_ram_56(0), A2 => gl_ram_n_823, B1 => gl_ram_ram_59(0), B2 => gl_ram_n_817, ZN => gl_ram_n_873);
  gl_ram_g13987 : AOI22D0BWP7T port map(A1 => gl_ram_ram_84(1), A2 => gl_ram_n_819, B1 => gl_ram_ram_85(1), B2 => gl_ram_n_818, ZN => gl_ram_n_872);
  gl_ram_g13988 : AOI22D0BWP7T port map(A1 => gl_ram_ram_54(0), A2 => gl_ram_n_826, B1 => gl_ram_ram_55(0), B2 => gl_ram_n_820, ZN => gl_ram_n_871);
  gl_ram_g13989 : AOI22D0BWP7T port map(A1 => gl_ram_ram_49(0), A2 => gl_ram_n_821, B1 => gl_ram_ram_50(0), B2 => gl_ram_n_825, ZN => gl_ram_n_870);
  gl_ram_g13990 : AOI22D0BWP7T port map(A1 => gl_ram_ram_80(1), A2 => gl_ram_n_823, B1 => gl_ram_ram_83(1), B2 => gl_ram_n_817, ZN => gl_ram_n_869);
  gl_ram_g13991 : AOI22D0BWP7T port map(A1 => gl_ram_ram_56(2), A2 => gl_ram_n_823, B1 => gl_ram_ram_59(2), B2 => gl_ram_n_817, ZN => gl_ram_n_868);
  gl_ram_g13992 : AOI22D0BWP7T port map(A1 => gl_ram_ram_52(0), A2 => gl_ram_n_819, B1 => gl_ram_ram_53(0), B2 => gl_ram_n_818, ZN => gl_ram_n_867);
  gl_ram_g13993 : AOI22D0BWP7T port map(A1 => gl_ram_ram_48(0), A2 => gl_ram_n_823, B1 => gl_ram_ram_51(0), B2 => gl_ram_n_817, ZN => gl_ram_n_866);
  gl_ram_g13994 : AOI22D0BWP7T port map(A1 => gl_ram_ram_81(2), A2 => gl_ram_n_821, B1 => gl_ram_ram_82(2), B2 => gl_ram_n_825, ZN => gl_ram_n_865);
  gl_ram_g13995 : AOI22D0BWP7T port map(A1 => gl_ram_ram_46(0), A2 => gl_ram_n_826, B1 => gl_ram_ram_47(0), B2 => gl_ram_n_820, ZN => gl_ram_n_864);
  gl_ram_g13996 : AOI22D0BWP7T port map(A1 => gl_ram_ram_78(1), A2 => gl_ram_n_826, B1 => gl_ram_ram_79(1), B2 => gl_ram_n_820, ZN => gl_ram_n_863);
  gl_ram_g13997 : AOI22D0BWP7T port map(A1 => gl_ram_ram_41(0), A2 => gl_ram_n_821, B1 => gl_ram_ram_42(0), B2 => gl_ram_n_825, ZN => gl_ram_n_862);
  gl_ram_g13998 : AOI22D0BWP7T port map(A1 => gl_ram_ram_72(1), A2 => gl_ram_n_823, B1 => gl_ram_ram_75(1), B2 => gl_ram_n_817, ZN => gl_ram_n_861);
  gl_ram_g13999 : AOI22D0BWP7T port map(A1 => gl_ram_ram_44(0), A2 => gl_ram_n_819, B1 => gl_ram_ram_45(0), B2 => gl_ram_n_818, ZN => gl_ram_n_860);
  gl_ram_g14000 : AOI22D0BWP7T port map(A1 => gl_ram_ram_40(0), A2 => gl_ram_n_823, B1 => gl_ram_ram_43(0), B2 => gl_ram_n_817, ZN => gl_ram_n_859);
  gl_ram_g14001 : AOI22D0BWP7T port map(A1 => gl_ram_ram_54(2), A2 => gl_ram_n_826, B1 => gl_ram_ram_55(2), B2 => gl_ram_n_820, ZN => gl_ram_n_858);
  gl_ram_g14002 : AOI22D0BWP7T port map(A1 => gl_ram_ram_76(1), A2 => gl_ram_n_819, B1 => gl_ram_ram_77(1), B2 => gl_ram_n_818, ZN => gl_ram_n_857);
  gl_ram_g14003 : AOI22D0BWP7T port map(A1 => gl_ram_ram_38(0), A2 => gl_ram_n_826, B1 => gl_ram_ram_39(0), B2 => gl_ram_n_820, ZN => gl_ram_n_856);
  gl_ram_g14004 : AOI22D0BWP7T port map(A1 => gl_ram_ram_73(1), A2 => gl_ram_n_821, B1 => gl_ram_ram_74(1), B2 => gl_ram_n_825, ZN => gl_ram_n_855);
  gl_ram_g14005 : AOI22D0BWP7T port map(A1 => gl_ram_ram_33(0), A2 => gl_ram_n_821, B1 => gl_ram_ram_34(0), B2 => gl_ram_n_825, ZN => gl_ram_n_854);
  gl_ram_g14006 : AOI22D0BWP7T port map(A1 => gl_ram_ram_36(0), A2 => gl_ram_n_819, B1 => gl_ram_ram_37(0), B2 => gl_ram_n_818, ZN => gl_ram_n_853);
  gl_ram_g14007 : AOI22D0BWP7T port map(A1 => gl_ram_ram_32(0), A2 => gl_ram_n_823, B1 => gl_ram_ram_35(0), B2 => gl_ram_n_817, ZN => gl_ram_n_852);
  gl_ram_g14008 : AOI22D0BWP7T port map(A1 => gl_ram_ram_48(2), A2 => gl_ram_n_823, B1 => gl_ram_ram_51(2), B2 => gl_ram_n_817, ZN => gl_ram_n_851);
  gl_ram_g14009 : AOI22D0BWP7T port map(A1 => gl_ram_ram_94(1), A2 => gl_ram_n_826, B1 => gl_ram_ram_95(1), B2 => gl_ram_n_820, ZN => gl_ram_n_850);
  gl_ram_g14010 : AOI22D0BWP7T port map(A1 => gl_ram_ram_30(0), A2 => gl_ram_n_826, B1 => gl_ram_ram_31(0), B2 => gl_ram_n_820, ZN => gl_ram_n_849);
  gl_ram_g14011 : AOI22D0BWP7T port map(A1 => gl_ram_ram_28(0), A2 => gl_ram_n_819, B1 => gl_ram_ram_29(0), B2 => gl_ram_n_818, ZN => gl_ram_n_848);
  gl_ram_g14012 : AOI22D0BWP7T port map(A1 => gl_ram_ram_89(1), A2 => gl_ram_n_821, B1 => gl_ram_ram_90(1), B2 => gl_ram_n_825, ZN => gl_ram_n_847);
  gl_ram_g14013 : AOI22D0BWP7T port map(A1 => gl_ram_ram_24(0), A2 => gl_ram_n_823, B1 => gl_ram_ram_27(0), B2 => gl_ram_n_817, ZN => gl_ram_n_846);
  gl_ram_g14014 : AOI22D0BWP7T port map(A1 => gl_ram_ram_52(2), A2 => gl_ram_n_819, B1 => gl_ram_ram_53(2), B2 => gl_ram_n_818, ZN => gl_ram_n_845);
  gl_ram_g14015 : AOI22D0BWP7T port map(A1 => gl_ram_ram_14(0), A2 => gl_ram_n_826, B1 => gl_ram_ram_15(0), B2 => gl_ram_n_820, ZN => gl_ram_n_844);
  gl_ram_g14016 : AOI22D0BWP7T port map(A1 => gl_ram_ram_8(0), A2 => gl_ram_n_823, B1 => gl_ram_ram_11(0), B2 => gl_ram_n_817, ZN => gl_ram_n_843);
  gl_ram_g14017 : AOI22D0BWP7T port map(A1 => gl_ram_ram_88(1), A2 => gl_ram_n_823, B1 => gl_ram_ram_91(1), B2 => gl_ram_n_817, ZN => gl_ram_n_842);
  gl_ram_g14018 : AOI22D0BWP7T port map(A1 => gl_ram_ram_12(0), A2 => gl_ram_n_819, B1 => gl_ram_ram_13(0), B2 => gl_ram_n_818, ZN => gl_ram_n_841);
  gl_ram_g14019 : AOI22D0BWP7T port map(A1 => gl_ram_ram_9(0), A2 => gl_ram_n_821, B1 => gl_ram_ram_10(0), B2 => gl_ram_n_825, ZN => gl_ram_n_840);
  gl_ram_g14020 : AOI22D0BWP7T port map(A1 => gl_ram_ram_70(1), A2 => gl_ram_n_826, B1 => gl_ram_ram_71(1), B2 => gl_ram_n_820, ZN => gl_ram_n_839);
  gl_ram_g14021 : AOI22D0BWP7T port map(A1 => gl_ram_ram_22(0), A2 => gl_ram_n_826, B1 => gl_ram_ram_23(0), B2 => gl_ram_n_820, ZN => gl_ram_n_838);
  gl_ram_g14022 : AOI22D0BWP7T port map(A1 => gl_ram_ram_20(0), A2 => gl_ram_n_819, B1 => gl_ram_ram_21(0), B2 => gl_ram_n_818, ZN => gl_ram_n_837);
  gl_ram_g14023 : AOI22D0BWP7T port map(A1 => gl_ram_ram_76(2), A2 => gl_ram_n_819, B1 => gl_ram_ram_77(2), B2 => gl_ram_n_818, ZN => gl_ram_n_836);
  gl_ram_g14024 : AOI22D0BWP7T port map(A1 => gl_ram_ram_68(1), A2 => gl_ram_n_819, B1 => gl_ram_ram_69(1), B2 => gl_ram_n_818, ZN => gl_ram_n_835);
  gl_ram_g14025 : AOI22D0BWP7T port map(A1 => gl_ram_ram_18(0), A2 => gl_ram_n_825, B1 => gl_ram_ram_19(0), B2 => gl_ram_n_817, ZN => gl_ram_n_834);
  gl_ram_g14026 : AOI22D0BWP7T port map(A1 => gl_ram_ram_16(0), A2 => gl_ram_n_823, B1 => gl_ram_ram_17(0), B2 => gl_ram_n_821, ZN => gl_ram_n_833);
  gl_ram_g14027 : AOI22D0BWP7T port map(A1 => gl_ram_ram_6(0), A2 => gl_ram_n_826, B1 => gl_ram_ram_7(0), B2 => gl_ram_n_820, ZN => gl_ram_n_832);
  gl_ram_g14028 : AOI22D0BWP7T port map(A1 => gl_ram_ram_46(2), A2 => gl_ram_n_826, B1 => gl_ram_ram_47(2), B2 => gl_ram_n_820, ZN => gl_ram_n_831);
  gl_ram_g14029 : AOI22D0BWP7T port map(A1 => gl_ram_ram_0(0), A2 => gl_ram_n_823, B1 => gl_ram_ram_3(0), B2 => gl_ram_n_817, ZN => gl_ram_n_830);
  gl_ram_g14030 : AOI22D0BWP7T port map(A1 => gl_ram_ram_4(0), A2 => gl_ram_n_819, B1 => gl_ram_ram_5(0), B2 => gl_ram_n_818, ZN => gl_ram_n_829);
  gl_ram_g14031 : AOI22D0BWP7T port map(A1 => gl_ram_ram_1(0), A2 => gl_ram_n_821, B1 => gl_ram_ram_2(0), B2 => gl_ram_n_825, ZN => gl_ram_n_828);
  gl_ram_g14032 : AOI22D0BWP7T port map(A1 => gl_ram_ram_6(2), A2 => gl_ram_n_826, B1 => gl_ram_ram_7(2), B2 => gl_ram_n_820, ZN => gl_ram_n_827);
  gl_ram_g14033 : INVD1BWP7T port map(I => gl_ram_n_824, ZN => gl_ram_n_825);
  gl_ram_g14034 : INVD1BWP7T port map(I => gl_ram_n_822, ZN => gl_ram_n_823);
  gl_ram_g14036 : AN2D1BWP7T port map(A1 => gl_ram_n_816, A2 => gl_ram_n_812, Z => gl_ram_n_826);
  gl_ram_g14037 : ND2D0BWP7T port map(A1 => gl_ram_n_815, A2 => gl_ram_n_812, ZN => gl_ram_n_824);
  gl_ram_g14038 : ND2D0BWP7T port map(A1 => gl_ram_n_815, A2 => gl_ram_n_810, ZN => gl_ram_n_822);
  gl_ram_g14039 : NR2XD0BWP7T port map(A1 => gl_ram_n_816, A2 => gl_ram_n_813, ZN => gl_ram_n_821);
  gl_ram_g14041 : NR2XD0BWP7T port map(A1 => gl_ram_n_815, A2 => gl_ram_n_811, ZN => gl_ram_n_820);
  gl_ram_g14042 : AN2D1BWP7T port map(A1 => gl_ram_n_816, A2 => gl_ram_n_810, Z => gl_ram_n_819);
  gl_ram_g14043 : NR2XD0BWP7T port map(A1 => gl_ram_n_815, A2 => gl_ram_n_813, ZN => gl_ram_n_818);
  gl_ram_g14044 : NR2XD0BWP7T port map(A1 => gl_ram_n_816, A2 => gl_ram_n_811, ZN => gl_ram_n_817);
  gl_ram_g14045 : INVD1BWP7T port map(I => gl_ram_n_816, ZN => gl_ram_n_815);
  gl_ram_g14046 : FA1D0BWP7T port map(A => gl_sig_x(2), B => gl_sig_y(1), CI => gl_ram_n_804, CO => gl_ram_n_814, S => gl_ram_n_816);
  gl_ram_g14047 : ND2D0BWP7T port map(A1 => gl_ram_n_805, A2 => gl_sig_x(0), ZN => gl_ram_n_813);
  gl_ram_g14048 : NR2D0BWP7T port map(A1 => gl_ram_n_805, A2 => gl_sig_x(0), ZN => gl_ram_n_812);
  gl_ram_g14049 : IND2D0BWP7T port map(A1 => gl_ram_n_805, B1 => gl_sig_x(0), ZN => gl_ram_n_811);
  gl_ram_g14050 : INR2D0BWP7T port map(A1 => gl_ram_n_805, B1 => gl_sig_x(0), ZN => gl_ram_n_810);
  gl_ram_g14051 : HA1D0BWP7T port map(A => gl_sig_x(3), B => gl_sig_y(0), CO => gl_ram_n_808, S => gl_ram_n_809);
  gl_ram_g14052 : HA1D0BWP7T port map(A => gl_sig_y(3), B => gl_sig_y(1), CO => gl_ram_n_806, S => gl_ram_n_807);
  gl_ram_g14053 : XNR2D1BWP7T port map(A1 => gl_sig_y(0), A2 => gl_sig_x(1), ZN => gl_ram_n_805);
  gl_ram_g14054 : AN2D1BWP7T port map(A1 => gl_sig_y(0), A2 => gl_sig_x(1), Z => gl_ram_n_804);
  gl_ram_g2 : INR2D1BWP7T port map(A1 => gl_ram_n_821, B1 => gl_ram_n_1023, ZN => gl_ram_n_803);
  gl_ram_g14055 : INR2D1BWP7T port map(A1 => gl_ram_n_817, B1 => gl_ram_n_1023, ZN => gl_ram_n_802);
  gl_ram_ram_position_reg_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_455, Q => gl_ram_ram_position(1));
  gl_ram_ram_position_reg_3 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_465, Q => gl_ram_ram_position(3));
  gl_ram_ram_position_reg_5 : DFQD0BWP7T port map(CP => clk, D => gl_ram_n_500, Q => gl_ram_ram_position(5));
  gl_ram_ram_position_reg_6 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_801, Q => gl_ram_ram_position(6));
  gl_ram_ram_reg_0_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_571, Q => gl_ram_ram_0(0));
  gl_ram_ram_reg_0_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_670, Q => gl_ram_ram_0(1));
  gl_ram_ram_reg_0_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_548, Q => gl_ram_ram_0(2));
  gl_ram_ram_reg_1_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_758, Q => gl_ram_ram_1(0));
  gl_ram_ram_reg_1_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_755, Q => gl_ram_ram_1(1));
  gl_ram_ram_reg_1_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_753, Q => gl_ram_ram_1(2));
  gl_ram_ram_reg_2_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_752, Q => gl_ram_ram_2(0));
  gl_ram_ram_reg_2_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_737, Q => gl_ram_ram_2(1));
  gl_ram_ram_reg_2_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_748, Q => gl_ram_ram_2(2));
  gl_ram_ram_reg_3_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_743, Q => gl_ram_ram_3(0));
  gl_ram_ram_reg_3_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_739, Q => gl_ram_ram_3(1));
  gl_ram_ram_reg_3_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_735, Q => gl_ram_ram_3(2));
  gl_ram_ram_reg_4_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_730, Q => gl_ram_ram_4(0));
  gl_ram_ram_reg_4_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_728, Q => gl_ram_ram_4(1));
  gl_ram_ram_reg_4_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_725, Q => gl_ram_ram_4(2));
  gl_ram_ram_reg_5_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_721, Q => gl_ram_ram_5(0));
  gl_ram_ram_reg_5_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_713, Q => gl_ram_ram_5(1));
  gl_ram_ram_reg_5_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_717, Q => gl_ram_ram_5(2));
  gl_ram_ram_reg_6_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_712, Q => gl_ram_ram_6(0));
  gl_ram_ram_reg_6_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_707, Q => gl_ram_ram_6(1));
  gl_ram_ram_reg_6_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_705, Q => gl_ram_ram_6(2));
  gl_ram_ram_reg_7_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_704, Q => gl_ram_ram_7(0));
  gl_ram_ram_reg_7_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_700, Q => gl_ram_ram_7(1));
  gl_ram_ram_reg_7_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_698, Q => gl_ram_ram_7(2));
  gl_ram_ram_reg_8_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_695, Q => gl_ram_ram_8(0));
  gl_ram_ram_reg_8_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_692, Q => gl_ram_ram_8(1));
  gl_ram_ram_reg_8_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_687, Q => gl_ram_ram_8(2));
  gl_ram_ram_reg_9_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_668, Q => gl_ram_ram_9(0));
  gl_ram_ram_reg_9_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_682, Q => gl_ram_ram_9(1));
  gl_ram_ram_reg_9_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_679, Q => gl_ram_ram_9(2));
  gl_ram_ram_reg_10_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_675, Q => gl_ram_ram_10(0));
  gl_ram_ram_reg_10_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_672, Q => gl_ram_ram_10(1));
  gl_ram_ram_reg_10_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_661, Q => gl_ram_ram_10(2));
  gl_ram_ram_reg_11_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_665, Q => gl_ram_ram_11(0));
  gl_ram_ram_reg_11_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_659, Q => gl_ram_ram_11(1));
  gl_ram_ram_reg_11_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_655, Q => gl_ram_ram_11(2));
  gl_ram_ram_reg_12_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_654, Q => gl_ram_ram_12(0));
  gl_ram_ram_reg_12_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_650, Q => gl_ram_ram_12(1));
  gl_ram_ram_reg_12_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_643, Q => gl_ram_ram_12(2));
  gl_ram_ram_reg_13_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_647, Q => gl_ram_ram_13(0));
  gl_ram_ram_reg_13_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_641, Q => gl_ram_ram_13(1));
  gl_ram_ram_reg_13_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_637, Q => gl_ram_ram_13(2));
  gl_ram_ram_reg_14_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_636, Q => gl_ram_ram_14(0));
  gl_ram_ram_reg_14_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_633, Q => gl_ram_ram_14(1));
  gl_ram_ram_reg_14_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_630, Q => gl_ram_ram_14(2));
  gl_ram_ram_reg_15_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_628, Q => gl_ram_ram_15(0));
  gl_ram_ram_reg_15_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_624, Q => gl_ram_ram_15(1));
  gl_ram_ram_reg_15_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_620, Q => gl_ram_ram_15(2));
  gl_ram_ram_reg_16_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_619, Q => gl_ram_ram_16(0));
  gl_ram_ram_reg_16_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_617, Q => gl_ram_ram_16(1));
  gl_ram_ram_reg_16_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_616, Q => gl_ram_ram_16(2));
  gl_ram_ram_reg_17_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_615, Q => gl_ram_ram_17(0));
  gl_ram_ram_reg_17_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_614, Q => gl_ram_ram_17(1));
  gl_ram_ram_reg_17_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_613, Q => gl_ram_ram_17(2));
  gl_ram_ram_reg_18_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_610, Q => gl_ram_ram_18(0));
  gl_ram_ram_reg_18_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_612, Q => gl_ram_ram_18(1));
  gl_ram_ram_reg_18_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_611, Q => gl_ram_ram_18(2));
  gl_ram_ram_reg_19_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_609, Q => gl_ram_ram_19(0));
  gl_ram_ram_reg_19_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_608, Q => gl_ram_ram_19(1));
  gl_ram_ram_reg_19_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_607, Q => gl_ram_ram_19(2));
  gl_ram_ram_reg_20_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_606, Q => gl_ram_ram_20(0));
  gl_ram_ram_reg_20_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_605, Q => gl_ram_ram_20(1));
  gl_ram_ram_reg_20_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_604, Q => gl_ram_ram_20(2));
  gl_ram_ram_reg_21_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_603, Q => gl_ram_ram_21(0));
  gl_ram_ram_reg_21_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_602, Q => gl_ram_ram_21(1));
  gl_ram_ram_reg_21_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_601, Q => gl_ram_ram_21(2));
  gl_ram_ram_reg_22_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_600, Q => gl_ram_ram_22(0));
  gl_ram_ram_reg_22_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_599, Q => gl_ram_ram_22(1));
  gl_ram_ram_reg_22_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_598, Q => gl_ram_ram_22(2));
  gl_ram_ram_reg_23_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_597, Q => gl_ram_ram_23(0));
  gl_ram_ram_reg_23_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_596, Q => gl_ram_ram_23(1));
  gl_ram_ram_reg_23_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_595, Q => gl_ram_ram_23(2));
  gl_ram_ram_reg_24_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_594, Q => gl_ram_ram_24(0));
  gl_ram_ram_reg_24_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_593, Q => gl_ram_ram_24(1));
  gl_ram_ram_reg_24_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_592, Q => gl_ram_ram_24(2));
  gl_ram_ram_reg_25_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_591, Q => gl_ram_ram_25(0));
  gl_ram_ram_reg_25_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_590, Q => gl_ram_ram_25(1));
  gl_ram_ram_reg_25_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_589, Q => gl_ram_ram_25(2));
  gl_ram_ram_reg_26_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_588, Q => gl_ram_ram_26(0));
  gl_ram_ram_reg_26_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_587, Q => gl_ram_ram_26(1));
  gl_ram_ram_reg_26_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_586, Q => gl_ram_ram_26(2));
  gl_ram_ram_reg_27_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_585, Q => gl_ram_ram_27(0));
  gl_ram_ram_reg_27_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_584, Q => gl_ram_ram_27(1));
  gl_ram_ram_reg_27_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_582, Q => gl_ram_ram_27(2));
  gl_ram_ram_reg_28_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_583, Q => gl_ram_ram_28(0));
  gl_ram_ram_reg_28_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_581, Q => gl_ram_ram_28(1));
  gl_ram_ram_reg_28_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_580, Q => gl_ram_ram_28(2));
  gl_ram_ram_reg_29_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_579, Q => gl_ram_ram_29(0));
  gl_ram_ram_reg_29_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_578, Q => gl_ram_ram_29(1));
  gl_ram_ram_reg_29_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_577, Q => gl_ram_ram_29(2));
  gl_ram_ram_reg_30_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_651, Q => gl_ram_ram_30(0));
  gl_ram_ram_reg_30_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_575, Q => gl_ram_ram_30(1));
  gl_ram_ram_reg_30_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_574, Q => gl_ram_ram_30(2));
  gl_ram_ram_reg_31_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_573, Q => gl_ram_ram_31(0));
  gl_ram_ram_reg_31_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_572, Q => gl_ram_ram_31(1));
  gl_ram_ram_reg_31_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_570, Q => gl_ram_ram_31(2));
  gl_ram_ram_reg_32_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_569, Q => gl_ram_ram_32(0));
  gl_ram_ram_reg_32_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_568, Q => gl_ram_ram_32(1));
  gl_ram_ram_reg_32_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_567, Q => gl_ram_ram_32(2));
  gl_ram_ram_reg_33_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_566, Q => gl_ram_ram_33(0));
  gl_ram_ram_reg_33_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_565, Q => gl_ram_ram_33(1));
  gl_ram_ram_reg_33_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_564, Q => gl_ram_ram_33(2));
  gl_ram_ram_reg_34_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_563, Q => gl_ram_ram_34(0));
  gl_ram_ram_reg_34_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_562, Q => gl_ram_ram_34(1));
  gl_ram_ram_reg_34_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_561, Q => gl_ram_ram_34(2));
  gl_ram_ram_reg_35_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_560, Q => gl_ram_ram_35(0));
  gl_ram_ram_reg_35_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_559, Q => gl_ram_ram_35(1));
  gl_ram_ram_reg_35_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_558, Q => gl_ram_ram_35(2));
  gl_ram_ram_reg_36_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_557, Q => gl_ram_ram_36(0));
  gl_ram_ram_reg_36_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_556, Q => gl_ram_ram_36(1));
  gl_ram_ram_reg_36_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_555, Q => gl_ram_ram_36(2));
  gl_ram_ram_reg_37_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_554, Q => gl_ram_ram_37(0));
  gl_ram_ram_reg_37_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_553, Q => gl_ram_ram_37(1));
  gl_ram_ram_reg_37_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_552, Q => gl_ram_ram_37(2));
  gl_ram_ram_reg_38_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_551, Q => gl_ram_ram_38(0));
  gl_ram_ram_reg_38_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_550, Q => gl_ram_ram_38(1));
  gl_ram_ram_reg_38_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_549, Q => gl_ram_ram_38(2));
  gl_ram_ram_reg_39_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_547, Q => gl_ram_ram_39(0));
  gl_ram_ram_reg_39_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_546, Q => gl_ram_ram_39(1));
  gl_ram_ram_reg_39_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_545, Q => gl_ram_ram_39(2));
  gl_ram_ram_reg_40_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_544, Q => gl_ram_ram_40(0));
  gl_ram_ram_reg_40_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_543, Q => gl_ram_ram_40(1));
  gl_ram_ram_reg_40_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_542, Q => gl_ram_ram_40(2));
  gl_ram_ram_reg_41_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_540, Q => gl_ram_ram_41(0));
  gl_ram_ram_reg_41_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_541, Q => gl_ram_ram_41(1));
  gl_ram_ram_reg_41_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_539, Q => gl_ram_ram_41(2));
  gl_ram_ram_reg_42_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_538, Q => gl_ram_ram_42(0));
  gl_ram_ram_reg_42_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_537, Q => gl_ram_ram_42(1));
  gl_ram_ram_reg_42_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_535, Q => gl_ram_ram_42(2));
  gl_ram_ram_reg_43_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_536, Q => gl_ram_ram_43(0));
  gl_ram_ram_reg_43_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_534, Q => gl_ram_ram_43(1));
  gl_ram_ram_reg_43_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_533, Q => gl_ram_ram_43(2));
  gl_ram_ram_reg_44_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_532, Q => gl_ram_ram_44(0));
  gl_ram_ram_reg_44_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_531, Q => gl_ram_ram_44(1));
  gl_ram_ram_reg_44_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_530, Q => gl_ram_ram_44(2));
  gl_ram_ram_reg_45_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_529, Q => gl_ram_ram_45(0));
  gl_ram_ram_reg_45_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_528, Q => gl_ram_ram_45(1));
  gl_ram_ram_reg_45_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_527, Q => gl_ram_ram_45(2));
  gl_ram_ram_reg_46_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_526, Q => gl_ram_ram_46(0));
  gl_ram_ram_reg_46_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_525, Q => gl_ram_ram_46(1));
  gl_ram_ram_reg_46_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_524, Q => gl_ram_ram_46(2));
  gl_ram_ram_reg_47_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_523, Q => gl_ram_ram_47(0));
  gl_ram_ram_reg_47_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_522, Q => gl_ram_ram_47(1));
  gl_ram_ram_reg_47_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_521, Q => gl_ram_ram_47(2));
  gl_ram_ram_reg_48_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_520, Q => gl_ram_ram_48(0));
  gl_ram_ram_reg_48_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_519, Q => gl_ram_ram_48(1));
  gl_ram_ram_reg_48_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_518, Q => gl_ram_ram_48(2));
  gl_ram_ram_reg_49_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_517, Q => gl_ram_ram_49(0));
  gl_ram_ram_reg_49_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_516, Q => gl_ram_ram_49(1));
  gl_ram_ram_reg_49_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_515, Q => gl_ram_ram_49(2));
  gl_ram_ram_reg_50_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_514, Q => gl_ram_ram_50(0));
  gl_ram_ram_reg_50_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_513, Q => gl_ram_ram_50(1));
  gl_ram_ram_reg_50_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_512, Q => gl_ram_ram_50(2));
  gl_ram_ram_reg_51_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_511, Q => gl_ram_ram_51(0));
  gl_ram_ram_reg_51_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_510, Q => gl_ram_ram_51(1));
  gl_ram_ram_reg_51_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_509, Q => gl_ram_ram_51(2));
  gl_ram_ram_reg_52_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_508, Q => gl_ram_ram_52(0));
  gl_ram_ram_reg_52_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_507, Q => gl_ram_ram_52(1));
  gl_ram_ram_reg_52_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_506, Q => gl_ram_ram_52(2));
  gl_ram_ram_reg_53_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_505, Q => gl_ram_ram_53(0));
  gl_ram_ram_reg_53_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_504, Q => gl_ram_ram_53(1));
  gl_ram_ram_reg_53_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_503, Q => gl_ram_ram_53(2));
  gl_ram_ram_reg_54_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_502, Q => gl_ram_ram_54(0));
  gl_ram_ram_reg_54_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_501, Q => gl_ram_ram_54(1));
  gl_ram_ram_reg_54_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_652, Q => gl_ram_ram_54(2));
  gl_ram_ram_reg_55_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_799, Q => gl_ram_ram_55(0));
  gl_ram_ram_reg_55_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_798, Q => gl_ram_ram_55(1));
  gl_ram_ram_reg_55_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_797, Q => gl_ram_ram_55(2));
  gl_ram_ram_reg_56_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_796, Q => gl_ram_ram_56(0));
  gl_ram_ram_reg_56_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_795, Q => gl_ram_ram_56(1));
  gl_ram_ram_reg_56_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_794, Q => gl_ram_ram_56(2));
  gl_ram_ram_reg_57_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_793, Q => gl_ram_ram_57(0));
  gl_ram_ram_reg_57_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_792, Q => gl_ram_ram_57(1));
  gl_ram_ram_reg_57_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_791, Q => gl_ram_ram_57(2));
  gl_ram_ram_reg_58_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_790, Q => gl_ram_ram_58(0));
  gl_ram_ram_reg_58_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_789, Q => gl_ram_ram_58(1));
  gl_ram_ram_reg_58_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_788, Q => gl_ram_ram_58(2));
  gl_ram_ram_reg_59_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_787, Q => gl_ram_ram_59(0));
  gl_ram_ram_reg_59_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_786, Q => gl_ram_ram_59(1));
  gl_ram_ram_reg_59_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_785, Q => gl_ram_ram_59(2));
  gl_ram_ram_reg_60_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_784, Q => gl_ram_ram_60(0));
  gl_ram_ram_reg_60_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_783, Q => gl_ram_ram_60(1));
  gl_ram_ram_reg_60_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_782, Q => gl_ram_ram_60(2));
  gl_ram_ram_reg_61_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_781, Q => gl_ram_ram_61(0));
  gl_ram_ram_reg_61_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_780, Q => gl_ram_ram_61(1));
  gl_ram_ram_reg_61_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_779, Q => gl_ram_ram_61(2));
  gl_ram_ram_reg_62_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_778, Q => gl_ram_ram_62(0));
  gl_ram_ram_reg_62_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_777, Q => gl_ram_ram_62(1));
  gl_ram_ram_reg_62_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_775, Q => gl_ram_ram_62(2));
  gl_ram_ram_reg_63_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_774, Q => gl_ram_ram_63(0));
  gl_ram_ram_reg_63_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_773, Q => gl_ram_ram_63(1));
  gl_ram_ram_reg_63_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_772, Q => gl_ram_ram_63(2));
  gl_ram_ram_reg_64_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_771, Q => gl_ram_ram_64(0));
  gl_ram_ram_reg_64_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_769, Q => gl_ram_ram_64(1));
  gl_ram_ram_reg_64_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_770, Q => gl_ram_ram_64(2));
  gl_ram_ram_reg_65_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_768, Q => gl_ram_ram_65(0));
  gl_ram_ram_reg_65_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_767, Q => gl_ram_ram_65(1));
  gl_ram_ram_reg_65_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_766, Q => gl_ram_ram_65(2));
  gl_ram_ram_reg_66_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_765, Q => gl_ram_ram_66(0));
  gl_ram_ram_reg_66_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_764, Q => gl_ram_ram_66(1));
  gl_ram_ram_reg_66_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_763, Q => gl_ram_ram_66(2));
  gl_ram_ram_reg_67_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_762, Q => gl_ram_ram_67(0));
  gl_ram_ram_reg_67_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_761, Q => gl_ram_ram_67(1));
  gl_ram_ram_reg_67_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_760, Q => gl_ram_ram_67(2));
  gl_ram_ram_reg_68_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_759, Q => gl_ram_ram_68(0));
  gl_ram_ram_reg_68_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_757, Q => gl_ram_ram_68(1));
  gl_ram_ram_reg_68_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_756, Q => gl_ram_ram_68(2));
  gl_ram_ram_reg_69_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_754, Q => gl_ram_ram_69(0));
  gl_ram_ram_reg_69_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_751, Q => gl_ram_ram_69(1));
  gl_ram_ram_reg_69_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_750, Q => gl_ram_ram_69(2));
  gl_ram_ram_reg_70_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_749, Q => gl_ram_ram_70(0));
  gl_ram_ram_reg_70_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_747, Q => gl_ram_ram_70(1));
  gl_ram_ram_reg_70_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_746, Q => gl_ram_ram_70(2));
  gl_ram_ram_reg_71_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_745, Q => gl_ram_ram_71(0));
  gl_ram_ram_reg_71_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_744, Q => gl_ram_ram_71(1));
  gl_ram_ram_reg_71_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_742, Q => gl_ram_ram_71(2));
  gl_ram_ram_reg_72_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_741, Q => gl_ram_ram_72(0));
  gl_ram_ram_reg_72_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_740, Q => gl_ram_ram_72(1));
  gl_ram_ram_reg_72_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_738, Q => gl_ram_ram_72(2));
  gl_ram_ram_reg_73_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_736, Q => gl_ram_ram_73(0));
  gl_ram_ram_reg_73_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_734, Q => gl_ram_ram_73(1));
  gl_ram_ram_reg_73_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_733, Q => gl_ram_ram_73(2));
  gl_ram_ram_reg_74_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_732, Q => gl_ram_ram_74(0));
  gl_ram_ram_reg_74_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_731, Q => gl_ram_ram_74(1));
  gl_ram_ram_reg_74_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_729, Q => gl_ram_ram_74(2));
  gl_ram_ram_reg_75_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_727, Q => gl_ram_ram_75(0));
  gl_ram_ram_reg_75_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_726, Q => gl_ram_ram_75(1));
  gl_ram_ram_reg_75_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_724, Q => gl_ram_ram_75(2));
  gl_ram_ram_reg_76_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_723, Q => gl_ram_ram_76(0));
  gl_ram_ram_reg_76_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_722, Q => gl_ram_ram_76(1));
  gl_ram_ram_reg_76_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_720, Q => gl_ram_ram_76(2));
  gl_ram_ram_reg_77_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_719, Q => gl_ram_ram_77(0));
  gl_ram_ram_reg_77_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_718, Q => gl_ram_ram_77(1));
  gl_ram_ram_reg_77_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_716, Q => gl_ram_ram_77(2));
  gl_ram_ram_reg_78_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_715, Q => gl_ram_ram_78(0));
  gl_ram_ram_reg_78_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_714, Q => gl_ram_ram_78(1));
  gl_ram_ram_reg_78_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_711, Q => gl_ram_ram_78(2));
  gl_ram_ram_reg_79_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_710, Q => gl_ram_ram_79(0));
  gl_ram_ram_reg_79_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_709, Q => gl_ram_ram_79(1));
  gl_ram_ram_reg_79_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_708, Q => gl_ram_ram_79(2));
  gl_ram_ram_reg_80_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_706, Q => gl_ram_ram_80(0));
  gl_ram_ram_reg_80_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_703, Q => gl_ram_ram_80(1));
  gl_ram_ram_reg_80_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_702, Q => gl_ram_ram_80(2));
  gl_ram_ram_reg_81_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_701, Q => gl_ram_ram_81(0));
  gl_ram_ram_reg_81_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_699, Q => gl_ram_ram_81(1));
  gl_ram_ram_reg_81_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_697, Q => gl_ram_ram_81(2));
  gl_ram_ram_reg_82_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_696, Q => gl_ram_ram_82(0));
  gl_ram_ram_reg_82_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_694, Q => gl_ram_ram_82(1));
  gl_ram_ram_reg_82_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_693, Q => gl_ram_ram_82(2));
  gl_ram_ram_reg_83_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_691, Q => gl_ram_ram_83(0));
  gl_ram_ram_reg_83_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_690, Q => gl_ram_ram_83(1));
  gl_ram_ram_reg_83_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_689, Q => gl_ram_ram_83(2));
  gl_ram_ram_reg_84_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_686, Q => gl_ram_ram_84(0));
  gl_ram_ram_reg_84_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_685, Q => gl_ram_ram_84(1));
  gl_ram_ram_reg_84_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_684, Q => gl_ram_ram_84(2));
  gl_ram_ram_reg_85_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_683, Q => gl_ram_ram_85(0));
  gl_ram_ram_reg_85_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_681, Q => gl_ram_ram_85(1));
  gl_ram_ram_reg_85_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_680, Q => gl_ram_ram_85(2));
  gl_ram_ram_reg_86_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_678, Q => gl_ram_ram_86(0));
  gl_ram_ram_reg_86_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_677, Q => gl_ram_ram_86(1));
  gl_ram_ram_reg_86_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_676, Q => gl_ram_ram_86(2));
  gl_ram_ram_reg_87_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_674, Q => gl_ram_ram_87(0));
  gl_ram_ram_reg_87_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_673, Q => gl_ram_ram_87(1));
  gl_ram_ram_reg_87_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_671, Q => gl_ram_ram_87(2));
  gl_ram_ram_reg_88_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_669, Q => gl_ram_ram_88(0));
  gl_ram_ram_reg_88_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_667, Q => gl_ram_ram_88(1));
  gl_ram_ram_reg_88_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_666, Q => gl_ram_ram_88(2));
  gl_ram_ram_reg_89_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_664, Q => gl_ram_ram_89(0));
  gl_ram_ram_reg_89_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_663, Q => gl_ram_ram_89(1));
  gl_ram_ram_reg_89_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_662, Q => gl_ram_ram_89(2));
  gl_ram_ram_reg_90_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_660, Q => gl_ram_ram_90(0));
  gl_ram_ram_reg_90_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_658, Q => gl_ram_ram_90(1));
  gl_ram_ram_reg_90_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_657, Q => gl_ram_ram_90(2));
  gl_ram_ram_reg_91_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_656, Q => gl_ram_ram_91(0));
  gl_ram_ram_reg_91_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_653, Q => gl_ram_ram_91(1));
  gl_ram_ram_reg_91_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_800, Q => gl_ram_ram_91(2));
  gl_ram_ram_reg_92_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_576, Q => gl_ram_ram_92(0));
  gl_ram_ram_reg_92_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_649, Q => gl_ram_ram_92(1));
  gl_ram_ram_reg_92_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_648, Q => gl_ram_ram_92(2));
  gl_ram_ram_reg_93_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_646, Q => gl_ram_ram_93(0));
  gl_ram_ram_reg_93_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_645, Q => gl_ram_ram_93(1));
  gl_ram_ram_reg_93_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_644, Q => gl_ram_ram_93(2));
  gl_ram_ram_reg_94_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_642, Q => gl_ram_ram_94(0));
  gl_ram_ram_reg_94_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_640, Q => gl_ram_ram_94(1));
  gl_ram_ram_reg_94_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_639, Q => gl_ram_ram_94(2));
  gl_ram_ram_reg_95_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_638, Q => gl_ram_ram_95(0));
  gl_ram_ram_reg_95_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_688, Q => gl_ram_ram_95(1));
  gl_ram_ram_reg_95_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_635, Q => gl_ram_ram_95(2));
  gl_ram_ram_reg_96_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_634, Q => gl_ram_ram_96(0));
  gl_ram_ram_reg_96_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_632, Q => gl_ram_ram_96(1));
  gl_ram_ram_reg_96_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_631, Q => gl_ram_ram_96(2));
  gl_ram_ram_reg_97_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_629, Q => gl_ram_ram_97(0));
  gl_ram_ram_reg_97_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_627, Q => gl_ram_ram_97(1));
  gl_ram_ram_reg_97_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_626, Q => gl_ram_ram_97(2));
  gl_ram_ram_reg_98_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_625, Q => gl_ram_ram_98(0));
  gl_ram_ram_reg_98_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_623, Q => gl_ram_ram_98(1));
  gl_ram_ram_reg_98_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_622, Q => gl_ram_ram_98(2));
  gl_ram_ram_reg_99_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_621, Q => gl_ram_ram_99(0));
  gl_ram_ram_reg_99_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_776, Q => gl_ram_ram_99(1));
  gl_ram_ram_reg_99_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_618, Q => gl_ram_ram_99(2));
  gl_ram_x_grid_reg_0 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_453, Q => gl_ram_x_grid(0));
  gl_ram_x_grid_reg_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_458, Q => gl_ram_x_grid(1));
  gl_ram_x_grid_reg_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_456, Q => gl_ram_x_grid(2));
  gl_ram_x_grid_reg_3 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_459, Q => gl_ram_x_grid(3));
  gl_ram_y_grid_reg_1 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_460, Q => gl_ram_y_grid(1));
  gl_ram_y_grid_reg_2 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_452, Q => gl_ram_y_grid(2));
  gl_ram_y_grid_reg_3 : DFQD1BWP7T port map(CP => clk, D => gl_ram_n_451, Q => gl_ram_y_grid(3));
  gl_ram_g27927 : MOAI22D0BWP7T port map(A1 => gl_ram_n_499, A2 => gl_ram_n_323, B1 => gl_ram_n_0, B2 => gl_ram_ram_position(6), ZN => gl_ram_n_801);
  gl_ram_g28078 : AO221D0BWP7T port map(A1 => gl_ram_n_484, A2 => gl_ram_n_273, B1 => gl_ram_n_446, B2 => gl_ram_ram_91(2), C => n_0, Z => gl_ram_n_800);
  gl_ram_g28079 : AO221D0BWP7T port map(A1 => gl_ram_n_489, A2 => gl_ram_n_282, B1 => gl_ram_n_410, B2 => gl_ram_ram_55(0), C => n_0, Z => gl_ram_n_799);
  gl_ram_g28080 : AO221D0BWP7T port map(A1 => gl_ram_n_490, A2 => gl_ram_n_282, B1 => gl_ram_n_410, B2 => gl_ram_ram_55(1), C => n_0, Z => gl_ram_n_798);
  gl_ram_g28081 : AO221D0BWP7T port map(A1 => gl_ram_n_491, A2 => gl_ram_n_282, B1 => gl_ram_n_410, B2 => gl_ram_ram_55(2), C => n_0, Z => gl_ram_n_797);
  gl_ram_g28082 : AO221D0BWP7T port map(A1 => gl_ram_n_473, A2 => gl_ram_n_287, B1 => gl_ram_n_413, B2 => gl_ram_ram_56(0), C => n_0, Z => gl_ram_n_796);
  gl_ram_g28083 : AO221D0BWP7T port map(A1 => gl_ram_n_492, A2 => gl_ram_n_287, B1 => gl_ram_n_413, B2 => gl_ram_ram_56(1), C => n_0, Z => gl_ram_n_795);
  gl_ram_g28084 : AO221D0BWP7T port map(A1 => gl_ram_n_474, A2 => gl_ram_n_287, B1 => gl_ram_n_413, B2 => gl_ram_ram_56(2), C => n_0, Z => gl_ram_n_794);
  gl_ram_g28085 : AO221D0BWP7T port map(A1 => gl_ram_n_473, A2 => gl_ram_n_285, B1 => gl_ram_n_409, B2 => gl_ram_ram_57(0), C => n_0, Z => gl_ram_n_793);
  gl_ram_g28086 : AO221D0BWP7T port map(A1 => gl_ram_n_492, A2 => gl_ram_n_285, B1 => gl_ram_n_409, B2 => gl_ram_ram_57(1), C => n_0, Z => gl_ram_n_792);
  gl_ram_g28087 : AO221D0BWP7T port map(A1 => gl_ram_n_474, A2 => gl_ram_n_285, B1 => gl_ram_n_409, B2 => gl_ram_ram_57(2), C => n_0, Z => gl_ram_n_791);
  gl_ram_g28088 : AO221D0BWP7T port map(A1 => gl_ram_n_473, A2 => gl_ram_n_286, B1 => gl_ram_n_352, B2 => gl_ram_ram_58(0), C => n_0, Z => gl_ram_n_790);
  gl_ram_g28089 : AO221D0BWP7T port map(A1 => gl_ram_n_492, A2 => gl_ram_n_286, B1 => gl_ram_n_352, B2 => gl_ram_ram_58(1), C => n_0, Z => gl_ram_n_789);
  gl_ram_g28090 : AO221D0BWP7T port map(A1 => gl_ram_n_474, A2 => gl_ram_n_286, B1 => gl_ram_n_352, B2 => gl_ram_ram_58(2), C => n_0, Z => gl_ram_n_788);
  gl_ram_g28091 : AO221D0BWP7T port map(A1 => gl_ram_n_473, A2 => gl_ram_n_284, B1 => gl_ram_n_408, B2 => gl_ram_ram_59(0), C => n_0, Z => gl_ram_n_787);
  gl_ram_g28092 : AO221D0BWP7T port map(A1 => gl_ram_n_492, A2 => gl_ram_n_284, B1 => gl_ram_n_408, B2 => gl_ram_ram_59(1), C => n_0, Z => gl_ram_n_786);
  gl_ram_g28093 : AO221D0BWP7T port map(A1 => gl_ram_n_474, A2 => gl_ram_n_284, B1 => gl_ram_n_408, B2 => gl_ram_ram_59(2), C => n_0, Z => gl_ram_n_785);
  gl_ram_g28094 : AO221D0BWP7T port map(A1 => gl_ram_n_489, A2 => gl_ram_n_287, B1 => gl_ram_n_407, B2 => gl_ram_ram_60(0), C => n_0, Z => gl_ram_n_784);
  gl_ram_g28095 : AO221D0BWP7T port map(A1 => gl_ram_n_490, A2 => gl_ram_n_287, B1 => gl_ram_n_407, B2 => gl_ram_ram_60(1), C => n_0, Z => gl_ram_n_783);
  gl_ram_g28096 : AO221D0BWP7T port map(A1 => gl_ram_n_491, A2 => gl_ram_n_287, B1 => gl_ram_n_407, B2 => gl_ram_ram_60(2), C => n_0, Z => gl_ram_n_782);
  gl_ram_g28097 : AO221D0BWP7T port map(A1 => gl_ram_n_489, A2 => gl_ram_n_285, B1 => gl_ram_n_405, B2 => gl_ram_ram_61(0), C => n_0, Z => gl_ram_n_781);
  gl_ram_g28098 : AO221D0BWP7T port map(A1 => gl_ram_n_490, A2 => gl_ram_n_285, B1 => gl_ram_n_405, B2 => gl_ram_ram_61(1), C => n_0, Z => gl_ram_n_780);
  gl_ram_g28099 : AO221D0BWP7T port map(A1 => gl_ram_n_491, A2 => gl_ram_n_285, B1 => gl_ram_n_405, B2 => gl_ram_ram_61(2), C => n_0, Z => gl_ram_n_779);
  gl_ram_g28100 : AO221D0BWP7T port map(A1 => gl_ram_n_489, A2 => gl_ram_n_286, B1 => gl_ram_n_356, B2 => gl_ram_ram_62(0), C => n_0, Z => gl_ram_n_778);
  gl_ram_g28101 : AO221D0BWP7T port map(A1 => gl_ram_n_490, A2 => gl_ram_n_286, B1 => gl_ram_n_356, B2 => gl_ram_ram_62(1), C => n_0, Z => gl_ram_n_777);
  gl_ram_g28102 : AO221D0BWP7T port map(A1 => gl_ram_n_480, A2 => gl_ram_n_282, B1 => gl_ram_n_372, B2 => gl_ram_ram_99(1), C => n_0, Z => gl_ram_n_776);
  gl_ram_g28103 : AO221D0BWP7T port map(A1 => gl_ram_n_491, A2 => gl_ram_n_286, B1 => gl_ram_n_356, B2 => gl_ram_ram_62(2), C => n_0, Z => gl_ram_n_775);
  gl_ram_g28104 : AO221D0BWP7T port map(A1 => gl_ram_n_489, A2 => gl_ram_n_284, B1 => gl_ram_n_406, B2 => gl_ram_ram_63(0), C => n_0, Z => gl_ram_n_774);
  gl_ram_g28105 : AO221D0BWP7T port map(A1 => gl_ram_n_490, A2 => gl_ram_n_284, B1 => gl_ram_n_406, B2 => gl_ram_ram_63(1), C => n_0, Z => gl_ram_n_773);
  gl_ram_g28106 : AO221D0BWP7T port map(A1 => gl_ram_n_491, A2 => gl_ram_n_284, B1 => gl_ram_n_406, B2 => gl_ram_ram_63(2), C => n_0, Z => gl_ram_n_772);
  gl_ram_g28107 : AO221D0BWP7T port map(A1 => gl_ram_n_479, A2 => gl_ram_n_277, B1 => gl_ram_n_428, B2 => gl_ram_ram_64(0), C => n_0, Z => gl_ram_n_771);
  gl_ram_g28108 : AO221D0BWP7T port map(A1 => gl_ram_n_481, A2 => gl_ram_n_277, B1 => gl_ram_n_428, B2 => gl_ram_ram_64(2), C => n_0, Z => gl_ram_n_770);
  gl_ram_g28109 : AO221D0BWP7T port map(A1 => gl_ram_n_480, A2 => gl_ram_n_277, B1 => gl_ram_n_428, B2 => gl_ram_ram_64(1), C => n_0, Z => gl_ram_n_769);
  gl_ram_g28110 : AO221D0BWP7T port map(A1 => gl_ram_n_479, A2 => gl_ram_n_274, B1 => gl_ram_n_368, B2 => gl_ram_ram_65(0), C => n_0, Z => gl_ram_n_768);
  gl_ram_g28111 : AO221D0BWP7T port map(A1 => gl_ram_n_480, A2 => gl_ram_n_274, B1 => gl_ram_n_368, B2 => gl_ram_ram_65(1), C => n_0, Z => gl_ram_n_767);
  gl_ram_g28112 : AO221D0BWP7T port map(A1 => gl_ram_n_481, A2 => gl_ram_n_274, B1 => gl_ram_n_368, B2 => gl_ram_ram_65(2), C => n_0, Z => gl_ram_n_766);
  gl_ram_g28113 : AO221D0BWP7T port map(A1 => gl_ram_n_479, A2 => gl_ram_n_275, B1 => gl_ram_n_418, B2 => gl_ram_ram_66(0), C => n_0, Z => gl_ram_n_765);
  gl_ram_g28114 : AO221D0BWP7T port map(A1 => gl_ram_n_480, A2 => gl_ram_n_275, B1 => gl_ram_n_418, B2 => gl_ram_ram_66(1), C => n_0, Z => gl_ram_n_764);
  gl_ram_g28115 : AO221D0BWP7T port map(A1 => gl_ram_n_481, A2 => gl_ram_n_275, B1 => gl_ram_n_418, B2 => gl_ram_ram_66(2), C => n_0, Z => gl_ram_n_763);
  gl_ram_g28116 : AO221D0BWP7T port map(A1 => gl_ram_n_479, A2 => gl_ram_n_276, B1 => gl_ram_n_361, B2 => gl_ram_ram_67(0), C => n_0, Z => gl_ram_n_762);
  gl_ram_g28117 : AO221D0BWP7T port map(A1 => gl_ram_n_480, A2 => gl_ram_n_276, B1 => gl_ram_n_361, B2 => gl_ram_ram_67(1), C => n_0, Z => gl_ram_n_761);
  gl_ram_g28118 : AO221D0BWP7T port map(A1 => gl_ram_n_481, A2 => gl_ram_n_276, B1 => gl_ram_n_361, B2 => gl_ram_ram_67(2), C => n_0, Z => gl_ram_n_760);
  gl_ram_g28119 : AO221D0BWP7T port map(A1 => gl_ram_n_482, A2 => gl_ram_n_277, B1 => gl_ram_n_444, B2 => gl_ram_ram_68(0), C => n_0, Z => gl_ram_n_759);
  gl_ram_g28120 : AO221D0BWP7T port map(A1 => gl_ram_n_476, A2 => gl_ram_n_274, B1 => gl_ram_n_359, B2 => gl_ram_ram_1(0), C => n_0, Z => gl_ram_n_758);
  gl_ram_g28121 : AO221D0BWP7T port map(A1 => gl_ram_n_497, A2 => gl_ram_n_277, B1 => gl_ram_n_444, B2 => gl_ram_ram_68(1), C => n_0, Z => gl_ram_n_757);
  gl_ram_g28122 : AO221D0BWP7T port map(A1 => gl_ram_n_483, A2 => gl_ram_n_277, B1 => gl_ram_n_444, B2 => gl_ram_ram_68(2), C => n_0, Z => gl_ram_n_756);
  gl_ram_g28123 : AO221D0BWP7T port map(A1 => gl_ram_n_488, A2 => gl_ram_n_274, B1 => gl_ram_n_359, B2 => gl_ram_ram_1(1), C => n_0, Z => gl_ram_n_755);
  gl_ram_g28124 : AO221D0BWP7T port map(A1 => gl_ram_n_482, A2 => gl_ram_n_274, B1 => gl_ram_n_450, B2 => gl_ram_ram_69(0), C => n_0, Z => gl_ram_n_754);
  gl_ram_g28125 : AO221D0BWP7T port map(A1 => gl_ram_n_475, A2 => gl_ram_n_274, B1 => gl_ram_n_359, B2 => gl_ram_ram_1(2), C => n_0, Z => gl_ram_n_753);
  gl_ram_g28126 : AO221D0BWP7T port map(A1 => gl_ram_n_476, A2 => gl_ram_n_275, B1 => gl_ram_n_390, B2 => gl_ram_ram_2(0), C => n_0, Z => gl_ram_n_752);
  gl_ram_g28127 : AO221D0BWP7T port map(A1 => gl_ram_n_497, A2 => gl_ram_n_274, B1 => gl_ram_n_450, B2 => gl_ram_ram_69(1), C => n_0, Z => gl_ram_n_751);
  gl_ram_g28128 : AO221D0BWP7T port map(A1 => gl_ram_n_483, A2 => gl_ram_n_274, B1 => gl_ram_n_450, B2 => gl_ram_ram_69(2), C => n_0, Z => gl_ram_n_750);
  gl_ram_g28129 : AO221D0BWP7T port map(A1 => gl_ram_n_482, A2 => gl_ram_n_275, B1 => gl_ram_n_440, B2 => gl_ram_ram_70(0), C => n_0, Z => gl_ram_n_749);
  gl_ram_g28130 : AO221D0BWP7T port map(A1 => gl_ram_n_475, A2 => gl_ram_n_275, B1 => gl_ram_n_390, B2 => gl_ram_ram_2(2), C => n_0, Z => gl_ram_n_748);
  gl_ram_g28131 : AO221D0BWP7T port map(A1 => gl_ram_n_497, A2 => gl_ram_n_275, B1 => gl_ram_n_440, B2 => gl_ram_ram_70(1), C => n_0, Z => gl_ram_n_747);
  gl_ram_g28132 : AO221D0BWP7T port map(A1 => gl_ram_n_483, A2 => gl_ram_n_275, B1 => gl_ram_n_440, B2 => gl_ram_ram_70(2), C => n_0, Z => gl_ram_n_746);
  gl_ram_g28133 : AO221D0BWP7T port map(A1 => gl_ram_n_482, A2 => gl_ram_n_276, B1 => gl_ram_n_434, B2 => gl_ram_ram_71(0), C => n_0, Z => gl_ram_n_745);
  gl_ram_g28134 : AO221D0BWP7T port map(A1 => gl_ram_n_497, A2 => gl_ram_n_276, B1 => gl_ram_n_434, B2 => gl_ram_ram_71(1), C => n_0, Z => gl_ram_n_744);
  gl_ram_g28135 : AO221D0BWP7T port map(A1 => gl_ram_n_476, A2 => gl_ram_n_276, B1 => gl_ram_n_377, B2 => gl_ram_ram_3(0), C => n_0, Z => gl_ram_n_743);
  gl_ram_g28136 : AO221D0BWP7T port map(A1 => gl_ram_n_483, A2 => gl_ram_n_276, B1 => gl_ram_n_434, B2 => gl_ram_ram_71(2), C => n_0, Z => gl_ram_n_742);
  gl_ram_g28137 : AO221D0BWP7T port map(A1 => gl_ram_n_479, A2 => gl_ram_n_278, B1 => gl_ram_n_416, B2 => gl_ram_ram_72(0), C => n_0, Z => gl_ram_n_741);
  gl_ram_g28138 : AO221D0BWP7T port map(A1 => gl_ram_n_480, A2 => gl_ram_n_278, B1 => gl_ram_n_416, B2 => gl_ram_ram_72(1), C => n_0, Z => gl_ram_n_740);
  gl_ram_g28139 : AO221D0BWP7T port map(A1 => gl_ram_n_488, A2 => gl_ram_n_276, B1 => gl_ram_n_377, B2 => gl_ram_ram_3(1), C => n_0, Z => gl_ram_n_739);
  gl_ram_g28140 : AO221D0BWP7T port map(A1 => gl_ram_n_481, A2 => gl_ram_n_278, B1 => gl_ram_n_416, B2 => gl_ram_ram_72(2), C => n_0, Z => gl_ram_n_738);
  gl_ram_g28141 : AO221D0BWP7T port map(A1 => gl_ram_n_488, A2 => gl_ram_n_275, B1 => gl_ram_n_390, B2 => gl_ram_ram_2(1), C => n_0, Z => gl_ram_n_737);
  gl_ram_g28142 : AO221D0BWP7T port map(A1 => gl_ram_n_479, A2 => gl_ram_n_272, B1 => gl_ram_n_353, B2 => gl_ram_ram_73(0), C => n_0, Z => gl_ram_n_736);
  gl_ram_g28143 : AO221D0BWP7T port map(A1 => gl_ram_n_475, A2 => gl_ram_n_276, B1 => gl_ram_n_377, B2 => gl_ram_ram_3(2), C => n_0, Z => gl_ram_n_735);
  gl_ram_g28144 : AO221D0BWP7T port map(A1 => gl_ram_n_480, A2 => gl_ram_n_272, B1 => gl_ram_n_353, B2 => gl_ram_ram_73(1), C => n_0, Z => gl_ram_n_734);
  gl_ram_g28145 : AO221D0BWP7T port map(A1 => gl_ram_n_481, A2 => gl_ram_n_272, B1 => gl_ram_n_353, B2 => gl_ram_ram_73(2), C => n_0, Z => gl_ram_n_733);
  gl_ram_g28146 : AO221D0BWP7T port map(A1 => gl_ram_n_479, A2 => gl_ram_n_279, B1 => gl_ram_n_417, B2 => gl_ram_ram_74(0), C => n_0, Z => gl_ram_n_732);
  gl_ram_g28147 : AO221D0BWP7T port map(A1 => gl_ram_n_480, A2 => gl_ram_n_279, B1 => gl_ram_n_417, B2 => gl_ram_ram_74(1), C => n_0, Z => gl_ram_n_731);
  gl_ram_g28148 : AO221D0BWP7T port map(A1 => gl_ram_n_478, A2 => gl_ram_n_277, B1 => gl_ram_n_383, B2 => gl_ram_ram_4(0), C => n_0, Z => gl_ram_n_730);
  gl_ram_g28149 : AO221D0BWP7T port map(A1 => gl_ram_n_481, A2 => gl_ram_n_279, B1 => gl_ram_n_417, B2 => gl_ram_ram_74(2), C => n_0, Z => gl_ram_n_729);
  gl_ram_g28150 : AO221D0BWP7T port map(A1 => gl_ram_n_493, A2 => gl_ram_n_277, B1 => gl_ram_n_383, B2 => gl_ram_ram_4(1), C => n_0, Z => gl_ram_n_728);
  gl_ram_g28151 : AO221D0BWP7T port map(A1 => gl_ram_n_479, A2 => gl_ram_n_273, B1 => gl_ram_n_375, B2 => gl_ram_ram_75(0), C => n_0, Z => gl_ram_n_727);
  gl_ram_g28152 : AO221D0BWP7T port map(A1 => gl_ram_n_480, A2 => gl_ram_n_273, B1 => gl_ram_n_375, B2 => gl_ram_ram_75(1), C => n_0, Z => gl_ram_n_726);
  gl_ram_g28153 : AO221D0BWP7T port map(A1 => gl_ram_n_477, A2 => gl_ram_n_277, B1 => gl_ram_n_383, B2 => gl_ram_ram_4(2), C => n_0, Z => gl_ram_n_725);
  gl_ram_g28154 : AO221D0BWP7T port map(A1 => gl_ram_n_481, A2 => gl_ram_n_273, B1 => gl_ram_n_375, B2 => gl_ram_ram_75(2), C => n_0, Z => gl_ram_n_724);
  gl_ram_g28155 : AO221D0BWP7T port map(A1 => gl_ram_n_482, A2 => gl_ram_n_278, B1 => gl_ram_n_437, B2 => gl_ram_ram_76(0), C => n_0, Z => gl_ram_n_723);
  gl_ram_g28156 : AO221D0BWP7T port map(A1 => gl_ram_n_497, A2 => gl_ram_n_278, B1 => gl_ram_n_437, B2 => gl_ram_ram_76(1), C => n_0, Z => gl_ram_n_722);
  gl_ram_g28157 : AO221D0BWP7T port map(A1 => gl_ram_n_478, A2 => gl_ram_n_274, B1 => gl_ram_n_381, B2 => gl_ram_ram_5(0), C => n_0, Z => gl_ram_n_721);
  gl_ram_g28158 : AO221D0BWP7T port map(A1 => gl_ram_n_483, A2 => gl_ram_n_278, B1 => gl_ram_n_437, B2 => gl_ram_ram_76(2), C => n_0, Z => gl_ram_n_720);
  gl_ram_g28159 : AO221D0BWP7T port map(A1 => gl_ram_n_482, A2 => gl_ram_n_272, B1 => gl_ram_n_426, B2 => gl_ram_ram_77(0), C => n_0, Z => gl_ram_n_719);
  gl_ram_g28160 : AO221D0BWP7T port map(A1 => gl_ram_n_497, A2 => gl_ram_n_272, B1 => gl_ram_n_426, B2 => gl_ram_ram_77(1), C => n_0, Z => gl_ram_n_718);
  gl_ram_g28161 : AO221D0BWP7T port map(A1 => gl_ram_n_477, A2 => gl_ram_n_274, B1 => gl_ram_n_381, B2 => gl_ram_ram_5(2), C => n_0, Z => gl_ram_n_717);
  gl_ram_g28162 : AO221D0BWP7T port map(A1 => gl_ram_n_483, A2 => gl_ram_n_272, B1 => gl_ram_n_426, B2 => gl_ram_ram_77(2), C => n_0, Z => gl_ram_n_716);
  gl_ram_g28163 : AO221D0BWP7T port map(A1 => gl_ram_n_482, A2 => gl_ram_n_279, B1 => gl_ram_n_439, B2 => gl_ram_ram_78(0), C => n_0, Z => gl_ram_n_715);
  gl_ram_g28164 : AO221D0BWP7T port map(A1 => gl_ram_n_497, A2 => gl_ram_n_279, B1 => gl_ram_n_439, B2 => gl_ram_ram_78(1), C => n_0, Z => gl_ram_n_714);
  gl_ram_g28165 : AO221D0BWP7T port map(A1 => gl_ram_n_493, A2 => gl_ram_n_274, B1 => gl_ram_n_381, B2 => gl_ram_ram_5(1), C => n_0, Z => gl_ram_n_713);
  gl_ram_g28166 : AO221D0BWP7T port map(A1 => gl_ram_n_478, A2 => gl_ram_n_275, B1 => gl_ram_n_371, B2 => gl_ram_ram_6(0), C => n_0, Z => gl_ram_n_712);
  gl_ram_g28167 : AO221D0BWP7T port map(A1 => gl_ram_n_483, A2 => gl_ram_n_279, B1 => gl_ram_n_439, B2 => gl_ram_ram_78(2), C => n_0, Z => gl_ram_n_711);
  gl_ram_g28168 : AO221D0BWP7T port map(A1 => gl_ram_n_482, A2 => gl_ram_n_273, B1 => gl_ram_n_442, B2 => gl_ram_ram_79(0), C => n_0, Z => gl_ram_n_710);
  gl_ram_g28169 : AO221D0BWP7T port map(A1 => gl_ram_n_497, A2 => gl_ram_n_273, B1 => gl_ram_n_442, B2 => gl_ram_ram_79(1), C => n_0, Z => gl_ram_n_709);
  gl_ram_g28170 : AO221D0BWP7T port map(A1 => gl_ram_n_483, A2 => gl_ram_n_273, B1 => gl_ram_n_442, B2 => gl_ram_ram_79(2), C => n_0, Z => gl_ram_n_708);
  gl_ram_g28171 : AO221D0BWP7T port map(A1 => gl_ram_n_493, A2 => gl_ram_n_275, B1 => gl_ram_n_371, B2 => gl_ram_ram_6(1), C => n_0, Z => gl_ram_n_707);
  gl_ram_g28172 : AO221D0BWP7T port map(A1 => gl_ram_n_485, A2 => gl_ram_n_277, B1 => gl_ram_n_433, B2 => gl_ram_ram_80(0), C => n_0, Z => gl_ram_n_706);
  gl_ram_g28173 : AO221D0BWP7T port map(A1 => gl_ram_n_477, A2 => gl_ram_n_275, B1 => gl_ram_n_371, B2 => gl_ram_ram_6(2), C => n_0, Z => gl_ram_n_705);
  gl_ram_g28174 : AO221D0BWP7T port map(A1 => gl_ram_n_478, A2 => gl_ram_n_276, B1 => gl_ram_n_395, B2 => gl_ram_ram_7(0), C => n_0, Z => gl_ram_n_704);
  gl_ram_g28175 : AO221D0BWP7T port map(A1 => gl_ram_n_498, A2 => gl_ram_n_277, B1 => gl_ram_n_433, B2 => gl_ram_ram_80(1), C => n_0, Z => gl_ram_n_703);
  gl_ram_g28176 : AO221D0BWP7T port map(A1 => gl_ram_n_484, A2 => gl_ram_n_277, B1 => gl_ram_n_433, B2 => gl_ram_ram_80(2), C => n_0, Z => gl_ram_n_702);
  gl_ram_g28177 : AO221D0BWP7T port map(A1 => gl_ram_n_485, A2 => gl_ram_n_274, B1 => gl_ram_n_438, B2 => gl_ram_ram_81(0), C => n_0, Z => gl_ram_n_701);
  gl_ram_g28178 : AO221D0BWP7T port map(A1 => gl_ram_n_493, A2 => gl_ram_n_276, B1 => gl_ram_n_395, B2 => gl_ram_ram_7(1), C => n_0, Z => gl_ram_n_700);
  gl_ram_g28179 : AO221D0BWP7T port map(A1 => gl_ram_n_498, A2 => gl_ram_n_274, B1 => gl_ram_n_438, B2 => gl_ram_ram_81(1), C => n_0, Z => gl_ram_n_699);
  gl_ram_g28180 : AO221D0BWP7T port map(A1 => gl_ram_n_477, A2 => gl_ram_n_276, B1 => gl_ram_n_395, B2 => gl_ram_ram_7(2), C => n_0, Z => gl_ram_n_698);
  gl_ram_g28181 : AO221D0BWP7T port map(A1 => gl_ram_n_484, A2 => gl_ram_n_274, B1 => gl_ram_n_438, B2 => gl_ram_ram_81(2), C => n_0, Z => gl_ram_n_697);
  gl_ram_g28182 : AO221D0BWP7T port map(A1 => gl_ram_n_485, A2 => gl_ram_n_275, B1 => gl_ram_n_427, B2 => gl_ram_ram_82(0), C => n_0, Z => gl_ram_n_696);
  gl_ram_g28183 : AO221D0BWP7T port map(A1 => gl_ram_n_476, A2 => gl_ram_n_278, B1 => gl_ram_n_392, B2 => gl_ram_ram_8(0), C => n_0, Z => gl_ram_n_695);
  gl_ram_g28184 : AO221D0BWP7T port map(A1 => gl_ram_n_498, A2 => gl_ram_n_275, B1 => gl_ram_n_427, B2 => gl_ram_ram_82(1), C => n_0, Z => gl_ram_n_694);
  gl_ram_g28185 : AO221D0BWP7T port map(A1 => gl_ram_n_484, A2 => gl_ram_n_275, B1 => gl_ram_n_427, B2 => gl_ram_ram_82(2), C => n_0, Z => gl_ram_n_693);
  gl_ram_g28186 : AO221D0BWP7T port map(A1 => gl_ram_n_488, A2 => gl_ram_n_278, B1 => gl_ram_n_392, B2 => gl_ram_ram_8(1), C => n_0, Z => gl_ram_n_692);
  gl_ram_g28187 : AO221D0BWP7T port map(A1 => gl_ram_n_485, A2 => gl_ram_n_276, B1 => gl_ram_n_445, B2 => gl_ram_ram_83(0), C => n_0, Z => gl_ram_n_691);
  gl_ram_g28188 : AO221D0BWP7T port map(A1 => gl_ram_n_498, A2 => gl_ram_n_276, B1 => gl_ram_n_445, B2 => gl_ram_ram_83(1), C => n_0, Z => gl_ram_n_690);
  gl_ram_g28189 : AO221D0BWP7T port map(A1 => gl_ram_n_484, A2 => gl_ram_n_276, B1 => gl_ram_n_445, B2 => gl_ram_ram_83(2), C => n_0, Z => gl_ram_n_689);
  gl_ram_g28190 : AO221D0BWP7T port map(A1 => gl_ram_n_496, A2 => gl_ram_n_273, B1 => gl_ram_n_423, B2 => gl_ram_ram_95(1), C => n_0, Z => gl_ram_n_688);
  gl_ram_g28191 : AO221D0BWP7T port map(A1 => gl_ram_n_475, A2 => gl_ram_n_278, B1 => gl_ram_n_392, B2 => gl_ram_ram_8(2), C => n_0, Z => gl_ram_n_687);
  gl_ram_g28192 : AO221D0BWP7T port map(A1 => gl_ram_n_495, A2 => gl_ram_n_277, B1 => gl_ram_n_366, B2 => gl_ram_ram_84(0), C => n_0, Z => gl_ram_n_686);
  gl_ram_g28193 : AO221D0BWP7T port map(A1 => gl_ram_n_496, A2 => gl_ram_n_277, B1 => gl_ram_n_366, B2 => gl_ram_ram_84(1), C => n_0, Z => gl_ram_n_685);
  gl_ram_g28194 : AO221D0BWP7T port map(A1 => gl_ram_n_494, A2 => gl_ram_n_277, B1 => gl_ram_n_366, B2 => gl_ram_ram_84(2), C => n_0, Z => gl_ram_n_684);
  gl_ram_g28195 : AO221D0BWP7T port map(A1 => gl_ram_n_495, A2 => gl_ram_n_274, B1 => gl_ram_n_449, B2 => gl_ram_ram_85(0), C => n_0, Z => gl_ram_n_683);
  gl_ram_g28196 : AO221D0BWP7T port map(A1 => gl_ram_n_488, A2 => gl_ram_n_272, B1 => gl_ram_n_358, B2 => gl_ram_ram_9(1), C => n_0, Z => gl_ram_n_682);
  gl_ram_g28197 : AO221D0BWP7T port map(A1 => gl_ram_n_496, A2 => gl_ram_n_274, B1 => gl_ram_n_449, B2 => gl_ram_ram_85(1), C => n_0, Z => gl_ram_n_681);
  gl_ram_g28198 : AO221D0BWP7T port map(A1 => gl_ram_n_494, A2 => gl_ram_n_274, B1 => gl_ram_n_449, B2 => gl_ram_ram_85(2), C => n_0, Z => gl_ram_n_680);
  gl_ram_g28199 : AO221D0BWP7T port map(A1 => gl_ram_n_475, A2 => gl_ram_n_272, B1 => gl_ram_n_358, B2 => gl_ram_ram_9(2), C => n_0, Z => gl_ram_n_679);
  gl_ram_g28200 : AO221D0BWP7T port map(A1 => gl_ram_n_495, A2 => gl_ram_n_275, B1 => gl_ram_n_382, B2 => gl_ram_ram_86(0), C => n_0, Z => gl_ram_n_678);
  gl_ram_g28201 : AO221D0BWP7T port map(A1 => gl_ram_n_496, A2 => gl_ram_n_275, B1 => gl_ram_n_382, B2 => gl_ram_ram_86(1), C => n_0, Z => gl_ram_n_677);
  gl_ram_g28202 : AO221D0BWP7T port map(A1 => gl_ram_n_494, A2 => gl_ram_n_275, B1 => gl_ram_n_382, B2 => gl_ram_ram_86(2), C => n_0, Z => gl_ram_n_676);
  gl_ram_g28203 : AO221D0BWP7T port map(A1 => gl_ram_n_476, A2 => gl_ram_n_279, B1 => gl_ram_n_391, B2 => gl_ram_ram_10(0), C => n_0, Z => gl_ram_n_675);
  gl_ram_g28204 : AO221D0BWP7T port map(A1 => gl_ram_n_495, A2 => gl_ram_n_276, B1 => gl_ram_n_447, B2 => gl_ram_ram_87(0), C => n_0, Z => gl_ram_n_674);
  gl_ram_g28205 : AO221D0BWP7T port map(A1 => gl_ram_n_496, A2 => gl_ram_n_276, B1 => gl_ram_n_447, B2 => gl_ram_ram_87(1), C => n_0, Z => gl_ram_n_673);
  gl_ram_g28206 : AO221D0BWP7T port map(A1 => gl_ram_n_488, A2 => gl_ram_n_279, B1 => gl_ram_n_391, B2 => gl_ram_ram_10(1), C => n_0, Z => gl_ram_n_672);
  gl_ram_g28207 : AO221D0BWP7T port map(A1 => gl_ram_n_494, A2 => gl_ram_n_276, B1 => gl_ram_n_447, B2 => gl_ram_ram_87(2), C => n_0, Z => gl_ram_n_671);
  gl_ram_g28208 : AO221D0BWP7T port map(A1 => gl_ram_n_488, A2 => gl_ram_n_277, B1 => gl_ram_n_414, B2 => gl_ram_ram_0(1), C => n_0, Z => gl_ram_n_670);
  gl_ram_g28209 : AO221D0BWP7T port map(A1 => gl_ram_n_485, A2 => gl_ram_n_278, B1 => gl_ram_n_424, B2 => gl_ram_ram_88(0), C => n_0, Z => gl_ram_n_669);
  gl_ram_g28210 : AO221D0BWP7T port map(A1 => gl_ram_n_476, A2 => gl_ram_n_272, B1 => gl_ram_n_358, B2 => gl_ram_ram_9(0), C => n_0, Z => gl_ram_n_668);
  gl_ram_g28211 : AO221D0BWP7T port map(A1 => gl_ram_n_498, A2 => gl_ram_n_278, B1 => gl_ram_n_424, B2 => gl_ram_ram_88(1), C => n_0, Z => gl_ram_n_667);
  gl_ram_g28212 : AO221D0BWP7T port map(A1 => gl_ram_n_484, A2 => gl_ram_n_278, B1 => gl_ram_n_424, B2 => gl_ram_ram_88(2), C => n_0, Z => gl_ram_n_666);
  gl_ram_g28213 : AO221D0BWP7T port map(A1 => gl_ram_n_476, A2 => gl_ram_n_273, B1 => gl_ram_n_388, B2 => gl_ram_ram_11(0), C => n_0, Z => gl_ram_n_665);
  gl_ram_g28214 : AO221D0BWP7T port map(A1 => gl_ram_n_485, A2 => gl_ram_n_272, B1 => gl_ram_n_436, B2 => gl_ram_ram_89(0), C => n_0, Z => gl_ram_n_664);
  gl_ram_g28215 : AO221D0BWP7T port map(A1 => gl_ram_n_498, A2 => gl_ram_n_272, B1 => gl_ram_n_436, B2 => gl_ram_ram_89(1), C => n_0, Z => gl_ram_n_663);
  gl_ram_g28216 : AO221D0BWP7T port map(A1 => gl_ram_n_484, A2 => gl_ram_n_272, B1 => gl_ram_n_436, B2 => gl_ram_ram_89(2), C => n_0, Z => gl_ram_n_662);
  gl_ram_g28217 : AO221D0BWP7T port map(A1 => gl_ram_n_475, A2 => gl_ram_n_279, B1 => gl_ram_n_391, B2 => gl_ram_ram_10(2), C => n_0, Z => gl_ram_n_661);
  gl_ram_g28218 : AO221D0BWP7T port map(A1 => gl_ram_n_485, A2 => gl_ram_n_279, B1 => gl_ram_n_425, B2 => gl_ram_ram_90(0), C => n_0, Z => gl_ram_n_660);
  gl_ram_g28219 : AO221D0BWP7T port map(A1 => gl_ram_n_488, A2 => gl_ram_n_273, B1 => gl_ram_n_388, B2 => gl_ram_ram_11(1), C => n_0, Z => gl_ram_n_659);
  gl_ram_g28220 : AO221D0BWP7T port map(A1 => gl_ram_n_498, A2 => gl_ram_n_279, B1 => gl_ram_n_425, B2 => gl_ram_ram_90(1), C => n_0, Z => gl_ram_n_658);
  gl_ram_g28221 : AO221D0BWP7T port map(A1 => gl_ram_n_484, A2 => gl_ram_n_279, B1 => gl_ram_n_425, B2 => gl_ram_ram_90(2), C => n_0, Z => gl_ram_n_657);
  gl_ram_g28222 : AO221D0BWP7T port map(A1 => gl_ram_n_485, A2 => gl_ram_n_273, B1 => gl_ram_n_446, B2 => gl_ram_ram_91(0), C => n_0, Z => gl_ram_n_656);
  gl_ram_g28223 : AO221D0BWP7T port map(A1 => gl_ram_n_475, A2 => gl_ram_n_273, B1 => gl_ram_n_388, B2 => gl_ram_ram_11(2), C => n_0, Z => gl_ram_n_655);
  gl_ram_g28224 : AO221D0BWP7T port map(A1 => gl_ram_n_478, A2 => gl_ram_n_278, B1 => gl_ram_n_370, B2 => gl_ram_ram_12(0), C => n_0, Z => gl_ram_n_654);
  gl_ram_g28225 : AO221D0BWP7T port map(A1 => gl_ram_n_498, A2 => gl_ram_n_273, B1 => gl_ram_n_446, B2 => gl_ram_ram_91(1), C => n_0, Z => gl_ram_n_653);
  gl_ram_g28226 : AO221D0BWP7T port map(A1 => gl_ram_n_491, A2 => gl_ram_n_280, B1 => gl_ram_n_363, B2 => gl_ram_ram_54(2), C => n_0, Z => gl_ram_n_652);
  gl_ram_g28228 : AO221D0BWP7T port map(A1 => gl_ram_n_489, A2 => gl_ram_n_279, B1 => gl_ram_n_384, B2 => gl_ram_ram_30(0), C => n_0, Z => gl_ram_n_651);
  gl_ram_g28229 : AO221D0BWP7T port map(A1 => gl_ram_n_493, A2 => gl_ram_n_278, B1 => gl_ram_n_370, B2 => gl_ram_ram_12(1), C => n_0, Z => gl_ram_n_650);
  gl_ram_g28230 : AO221D0BWP7T port map(A1 => gl_ram_n_496, A2 => gl_ram_n_278, B1 => gl_ram_n_365, B2 => gl_ram_ram_92(1), C => n_0, Z => gl_ram_n_649);
  gl_ram_g28231 : AO221D0BWP7T port map(A1 => gl_ram_n_494, A2 => gl_ram_n_278, B1 => gl_ram_n_365, B2 => gl_ram_ram_92(2), C => n_0, Z => gl_ram_n_648);
  gl_ram_g28232 : AO221D0BWP7T port map(A1 => gl_ram_n_478, A2 => gl_ram_n_272, B1 => gl_ram_n_380, B2 => gl_ram_ram_13(0), C => n_0, Z => gl_ram_n_647);
  gl_ram_g28233 : AO221D0BWP7T port map(A1 => gl_ram_n_495, A2 => gl_ram_n_272, B1 => gl_ram_n_448, B2 => gl_ram_ram_93(0), C => n_0, Z => gl_ram_n_646);
  gl_ram_g28234 : AO221D0BWP7T port map(A1 => gl_ram_n_496, A2 => gl_ram_n_272, B1 => gl_ram_n_448, B2 => gl_ram_ram_93(1), C => n_0, Z => gl_ram_n_645);
  gl_ram_g28235 : AO221D0BWP7T port map(A1 => gl_ram_n_494, A2 => gl_ram_n_272, B1 => gl_ram_n_448, B2 => gl_ram_ram_93(2), C => n_0, Z => gl_ram_n_644);
  gl_ram_g28236 : AO221D0BWP7T port map(A1 => gl_ram_n_477, A2 => gl_ram_n_278, B1 => gl_ram_n_370, B2 => gl_ram_ram_12(2), C => n_0, Z => gl_ram_n_643);
  gl_ram_g28237 : AO221D0BWP7T port map(A1 => gl_ram_n_495, A2 => gl_ram_n_279, B1 => gl_ram_n_411, B2 => gl_ram_ram_94(0), C => n_0, Z => gl_ram_n_642);
  gl_ram_g28238 : AO221D0BWP7T port map(A1 => gl_ram_n_493, A2 => gl_ram_n_272, B1 => gl_ram_n_380, B2 => gl_ram_ram_13(1), C => n_0, Z => gl_ram_n_641);
  gl_ram_g28239 : AO221D0BWP7T port map(A1 => gl_ram_n_496, A2 => gl_ram_n_279, B1 => gl_ram_n_411, B2 => gl_ram_ram_94(1), C => n_0, Z => gl_ram_n_640);
  gl_ram_g28240 : AO221D0BWP7T port map(A1 => gl_ram_n_494, A2 => gl_ram_n_279, B1 => gl_ram_n_411, B2 => gl_ram_ram_94(2), C => n_0, Z => gl_ram_n_639);
  gl_ram_g28241 : AO221D0BWP7T port map(A1 => gl_ram_n_495, A2 => gl_ram_n_273, B1 => gl_ram_n_423, B2 => gl_ram_ram_95(0), C => n_0, Z => gl_ram_n_638);
  gl_ram_g28242 : AO221D0BWP7T port map(A1 => gl_ram_n_477, A2 => gl_ram_n_272, B1 => gl_ram_n_380, B2 => gl_ram_ram_13(2), C => n_0, Z => gl_ram_n_637);
  gl_ram_g28243 : AO221D0BWP7T port map(A1 => gl_ram_n_478, A2 => gl_ram_n_279, B1 => gl_ram_n_374, B2 => gl_ram_ram_14(0), C => n_0, Z => gl_ram_n_636);
  gl_ram_g28244 : AO221D0BWP7T port map(A1 => gl_ram_n_494, A2 => gl_ram_n_273, B1 => gl_ram_n_423, B2 => gl_ram_ram_95(2), C => n_0, Z => gl_ram_n_635);
  gl_ram_g28245 : AO221D0BWP7T port map(A1 => gl_ram_n_479, A2 => gl_ram_n_281, B1 => gl_ram_n_443, B2 => gl_ram_ram_96(0), C => n_0, Z => gl_ram_n_634);
  gl_ram_g28246 : AO221D0BWP7T port map(A1 => gl_ram_n_493, A2 => gl_ram_n_279, B1 => gl_ram_n_374, B2 => gl_ram_ram_14(1), C => n_0, Z => gl_ram_n_633);
  gl_ram_g28247 : AO221D0BWP7T port map(A1 => gl_ram_n_480, A2 => gl_ram_n_281, B1 => gl_ram_n_443, B2 => gl_ram_ram_96(1), C => n_0, Z => gl_ram_n_632);
  gl_ram_g28248 : AO221D0BWP7T port map(A1 => gl_ram_n_481, A2 => gl_ram_n_281, B1 => gl_ram_n_443, B2 => gl_ram_ram_96(2), C => n_0, Z => gl_ram_n_631);
  gl_ram_g28249 : AO221D0BWP7T port map(A1 => gl_ram_n_477, A2 => gl_ram_n_279, B1 => gl_ram_n_374, B2 => gl_ram_ram_14(2), C => n_0, Z => gl_ram_n_630);
  gl_ram_g28250 : AO221D0BWP7T port map(A1 => gl_ram_n_479, A2 => gl_ram_n_283, B1 => gl_ram_n_412, B2 => gl_ram_ram_97(0), C => n_0, Z => gl_ram_n_629);
  gl_ram_g28251 : AO221D0BWP7T port map(A1 => gl_ram_n_478, A2 => gl_ram_n_273, B1 => gl_ram_n_415, B2 => gl_ram_ram_15(0), C => n_0, Z => gl_ram_n_628);
  gl_ram_g28252 : AO221D0BWP7T port map(A1 => gl_ram_n_480, A2 => gl_ram_n_283, B1 => gl_ram_n_412, B2 => gl_ram_ram_97(1), C => n_0, Z => gl_ram_n_627);
  gl_ram_g28253 : AO221D0BWP7T port map(A1 => gl_ram_n_481, A2 => gl_ram_n_283, B1 => gl_ram_n_412, B2 => gl_ram_ram_97(2), C => n_0, Z => gl_ram_n_626);
  gl_ram_g28254 : AO221D0BWP7T port map(A1 => gl_ram_n_479, A2 => gl_ram_n_280, B1 => gl_ram_n_432, B2 => gl_ram_ram_98(0), C => n_0, Z => gl_ram_n_625);
  gl_ram_g28255 : AO221D0BWP7T port map(A1 => gl_ram_n_493, A2 => gl_ram_n_273, B1 => gl_ram_n_415, B2 => gl_ram_ram_15(1), C => n_0, Z => gl_ram_n_624);
  gl_ram_g28256 : AO221D0BWP7T port map(A1 => gl_ram_n_480, A2 => gl_ram_n_280, B1 => gl_ram_n_432, B2 => gl_ram_ram_98(1), C => n_0, Z => gl_ram_n_623);
  gl_ram_g28257 : AO221D0BWP7T port map(A1 => gl_ram_n_481, A2 => gl_ram_n_280, B1 => gl_ram_n_432, B2 => gl_ram_ram_98(2), C => n_0, Z => gl_ram_n_622);
  gl_ram_g28258 : AO221D0BWP7T port map(A1 => gl_ram_n_479, A2 => gl_ram_n_282, B1 => gl_ram_n_372, B2 => gl_ram_ram_99(0), C => n_0, Z => gl_ram_n_621);
  gl_ram_g28259 : AO221D0BWP7T port map(A1 => gl_ram_n_477, A2 => gl_ram_n_273, B1 => gl_ram_n_415, B2 => gl_ram_ram_15(2), C => n_0, Z => gl_ram_n_620);
  gl_ram_g28260 : AO221D0BWP7T port map(A1 => gl_ram_n_473, A2 => gl_ram_n_277, B1 => gl_ram_n_362, B2 => gl_ram_ram_16(0), C => n_0, Z => gl_ram_n_619);
  gl_ram_g28261 : AO221D0BWP7T port map(A1 => gl_ram_n_481, A2 => gl_ram_n_282, B1 => gl_ram_n_372, B2 => gl_ram_ram_99(2), C => n_0, Z => gl_ram_n_618);
  gl_ram_g28262 : AO221D0BWP7T port map(A1 => gl_ram_n_492, A2 => gl_ram_n_277, B1 => gl_ram_n_362, B2 => gl_ram_ram_16(1), C => n_0, Z => gl_ram_n_617);
  gl_ram_g28263 : AO221D0BWP7T port map(A1 => gl_ram_n_474, A2 => gl_ram_n_277, B1 => gl_ram_n_362, B2 => gl_ram_ram_16(2), C => n_0, Z => gl_ram_n_616);
  gl_ram_g28264 : AO221D0BWP7T port map(A1 => gl_ram_n_473, A2 => gl_ram_n_274, B1 => gl_ram_n_404, B2 => gl_ram_ram_17(0), C => n_0, Z => gl_ram_n_615);
  gl_ram_g28265 : AO221D0BWP7T port map(A1 => gl_ram_n_492, A2 => gl_ram_n_274, B1 => gl_ram_n_404, B2 => gl_ram_ram_17(1), C => n_0, Z => gl_ram_n_614);
  gl_ram_g28266 : AO221D0BWP7T port map(A1 => gl_ram_n_474, A2 => gl_ram_n_274, B1 => gl_ram_n_404, B2 => gl_ram_ram_17(2), C => n_0, Z => gl_ram_n_613);
  gl_ram_g28267 : AO221D0BWP7T port map(A1 => gl_ram_n_492, A2 => gl_ram_n_275, B1 => gl_ram_n_360, B2 => gl_ram_ram_18(1), C => n_0, Z => gl_ram_n_612);
  gl_ram_g28268 : AO221D0BWP7T port map(A1 => gl_ram_n_474, A2 => gl_ram_n_275, B1 => gl_ram_n_360, B2 => gl_ram_ram_18(2), C => n_0, Z => gl_ram_n_611);
  gl_ram_g28269 : AO221D0BWP7T port map(A1 => gl_ram_n_473, A2 => gl_ram_n_275, B1 => gl_ram_n_360, B2 => gl_ram_ram_18(0), C => n_0, Z => gl_ram_n_610);
  gl_ram_g28270 : AO221D0BWP7T port map(A1 => gl_ram_n_473, A2 => gl_ram_n_276, B1 => gl_ram_n_421, B2 => gl_ram_ram_19(0), C => n_0, Z => gl_ram_n_609);
  gl_ram_g28271 : AO221D0BWP7T port map(A1 => gl_ram_n_492, A2 => gl_ram_n_276, B1 => gl_ram_n_421, B2 => gl_ram_ram_19(1), C => n_0, Z => gl_ram_n_608);
  gl_ram_g28272 : AO221D0BWP7T port map(A1 => gl_ram_n_474, A2 => gl_ram_n_276, B1 => gl_ram_n_421, B2 => gl_ram_ram_19(2), C => n_0, Z => gl_ram_n_607);
  gl_ram_g28273 : AO221D0BWP7T port map(A1 => gl_ram_n_489, A2 => gl_ram_n_277, B1 => gl_ram_n_355, B2 => gl_ram_ram_20(0), C => n_0, Z => gl_ram_n_606);
  gl_ram_g28274 : AO221D0BWP7T port map(A1 => gl_ram_n_490, A2 => gl_ram_n_277, B1 => gl_ram_n_355, B2 => gl_ram_ram_20(1), C => n_0, Z => gl_ram_n_605);
  gl_ram_g28275 : AO221D0BWP7T port map(A1 => gl_ram_n_491, A2 => gl_ram_n_277, B1 => gl_ram_n_355, B2 => gl_ram_ram_20(2), C => n_0, Z => gl_ram_n_604);
  gl_ram_g28276 : AO221D0BWP7T port map(A1 => gl_ram_n_489, A2 => gl_ram_n_274, B1 => gl_ram_n_403, B2 => gl_ram_ram_21(0), C => n_0, Z => gl_ram_n_603);
  gl_ram_g28277 : AO221D0BWP7T port map(A1 => gl_ram_n_490, A2 => gl_ram_n_274, B1 => gl_ram_n_403, B2 => gl_ram_ram_21(1), C => n_0, Z => gl_ram_n_602);
  gl_ram_g28278 : AO221D0BWP7T port map(A1 => gl_ram_n_491, A2 => gl_ram_n_274, B1 => gl_ram_n_403, B2 => gl_ram_ram_21(2), C => n_0, Z => gl_ram_n_601);
  gl_ram_g28279 : AO221D0BWP7T port map(A1 => gl_ram_n_489, A2 => gl_ram_n_275, B1 => gl_ram_n_376, B2 => gl_ram_ram_22(0), C => n_0, Z => gl_ram_n_600);
  gl_ram_g28280 : AO221D0BWP7T port map(A1 => gl_ram_n_490, A2 => gl_ram_n_275, B1 => gl_ram_n_376, B2 => gl_ram_ram_22(1), C => n_0, Z => gl_ram_n_599);
  gl_ram_g28281 : AO221D0BWP7T port map(A1 => gl_ram_n_491, A2 => gl_ram_n_275, B1 => gl_ram_n_376, B2 => gl_ram_ram_22(2), C => n_0, Z => gl_ram_n_598);
  gl_ram_g28282 : AO221D0BWP7T port map(A1 => gl_ram_n_489, A2 => gl_ram_n_276, B1 => gl_ram_n_420, B2 => gl_ram_ram_23(0), C => n_0, Z => gl_ram_n_597);
  gl_ram_g28283 : AO221D0BWP7T port map(A1 => gl_ram_n_490, A2 => gl_ram_n_276, B1 => gl_ram_n_420, B2 => gl_ram_ram_23(1), C => n_0, Z => gl_ram_n_596);
  gl_ram_g28284 : AO221D0BWP7T port map(A1 => gl_ram_n_491, A2 => gl_ram_n_276, B1 => gl_ram_n_420, B2 => gl_ram_ram_23(2), C => n_0, Z => gl_ram_n_595);
  gl_ram_g28285 : AO221D0BWP7T port map(A1 => gl_ram_n_473, A2 => gl_ram_n_278, B1 => gl_ram_n_351, B2 => gl_ram_ram_24(0), C => n_0, Z => gl_ram_n_594);
  gl_ram_g28286 : AO221D0BWP7T port map(A1 => gl_ram_n_492, A2 => gl_ram_n_278, B1 => gl_ram_n_351, B2 => gl_ram_ram_24(1), C => n_0, Z => gl_ram_n_593);
  gl_ram_g28287 : AO221D0BWP7T port map(A1 => gl_ram_n_474, A2 => gl_ram_n_278, B1 => gl_ram_n_351, B2 => gl_ram_ram_24(2), C => n_0, Z => gl_ram_n_592);
  gl_ram_g28288 : AO221D0BWP7T port map(A1 => gl_ram_n_473, A2 => gl_ram_n_272, B1 => gl_ram_n_402, B2 => gl_ram_ram_25(0), C => n_0, Z => gl_ram_n_591);
  gl_ram_g28289 : AO221D0BWP7T port map(A1 => gl_ram_n_492, A2 => gl_ram_n_272, B1 => gl_ram_n_402, B2 => gl_ram_ram_25(1), C => n_0, Z => gl_ram_n_590);
  gl_ram_g28290 : AO221D0BWP7T port map(A1 => gl_ram_n_474, A2 => gl_ram_n_272, B1 => gl_ram_n_402, B2 => gl_ram_ram_25(2), C => n_0, Z => gl_ram_n_589);
  gl_ram_g28291 : AO221D0BWP7T port map(A1 => gl_ram_n_473, A2 => gl_ram_n_279, B1 => gl_ram_n_373, B2 => gl_ram_ram_26(0), C => n_0, Z => gl_ram_n_588);
  gl_ram_g28292 : AO221D0BWP7T port map(A1 => gl_ram_n_492, A2 => gl_ram_n_279, B1 => gl_ram_n_373, B2 => gl_ram_ram_26(1), C => n_0, Z => gl_ram_n_587);
  gl_ram_g28293 : AO221D0BWP7T port map(A1 => gl_ram_n_474, A2 => gl_ram_n_279, B1 => gl_ram_n_373, B2 => gl_ram_ram_26(2), C => n_0, Z => gl_ram_n_586);
  gl_ram_g28294 : AO221D0BWP7T port map(A1 => gl_ram_n_473, A2 => gl_ram_n_273, B1 => gl_ram_n_431, B2 => gl_ram_ram_27(0), C => n_0, Z => gl_ram_n_585);
  gl_ram_g28295 : AO221D0BWP7T port map(A1 => gl_ram_n_492, A2 => gl_ram_n_273, B1 => gl_ram_n_431, B2 => gl_ram_ram_27(1), C => n_0, Z => gl_ram_n_584);
  gl_ram_g28296 : AO221D0BWP7T port map(A1 => gl_ram_n_489, A2 => gl_ram_n_278, B1 => gl_ram_n_354, B2 => gl_ram_ram_28(0), C => n_0, Z => gl_ram_n_583);
  gl_ram_g28297 : AO221D0BWP7T port map(A1 => gl_ram_n_474, A2 => gl_ram_n_273, B1 => gl_ram_n_431, B2 => gl_ram_ram_27(2), C => n_0, Z => gl_ram_n_582);
  gl_ram_g28298 : AO221D0BWP7T port map(A1 => gl_ram_n_490, A2 => gl_ram_n_278, B1 => gl_ram_n_354, B2 => gl_ram_ram_28(1), C => n_0, Z => gl_ram_n_581);
  gl_ram_g28299 : AO221D0BWP7T port map(A1 => gl_ram_n_491, A2 => gl_ram_n_278, B1 => gl_ram_n_354, B2 => gl_ram_ram_28(2), C => n_0, Z => gl_ram_n_580);
  gl_ram_g28300 : AO221D0BWP7T port map(A1 => gl_ram_n_489, A2 => gl_ram_n_272, B1 => gl_ram_n_400, B2 => gl_ram_ram_29(0), C => n_0, Z => gl_ram_n_579);
  gl_ram_g28301 : AO221D0BWP7T port map(A1 => gl_ram_n_490, A2 => gl_ram_n_272, B1 => gl_ram_n_400, B2 => gl_ram_ram_29(1), C => n_0, Z => gl_ram_n_578);
  gl_ram_g28302 : AO221D0BWP7T port map(A1 => gl_ram_n_491, A2 => gl_ram_n_272, B1 => gl_ram_n_400, B2 => gl_ram_ram_29(2), C => n_0, Z => gl_ram_n_577);
  gl_ram_g28303 : AO221D0BWP7T port map(A1 => gl_ram_n_495, A2 => gl_ram_n_278, B1 => gl_ram_n_365, B2 => gl_ram_ram_92(0), C => n_0, Z => gl_ram_n_576);
  gl_ram_g28304 : AO221D0BWP7T port map(A1 => gl_ram_n_490, A2 => gl_ram_n_279, B1 => gl_ram_n_384, B2 => gl_ram_ram_30(1), C => n_0, Z => gl_ram_n_575);
  gl_ram_g28305 : AO221D0BWP7T port map(A1 => gl_ram_n_491, A2 => gl_ram_n_279, B1 => gl_ram_n_384, B2 => gl_ram_ram_30(2), C => n_0, Z => gl_ram_n_574);
  gl_ram_g28306 : AO221D0BWP7T port map(A1 => gl_ram_n_489, A2 => gl_ram_n_273, B1 => gl_ram_n_430, B2 => gl_ram_ram_31(0), C => n_0, Z => gl_ram_n_573);
  gl_ram_g28307 : AO221D0BWP7T port map(A1 => gl_ram_n_490, A2 => gl_ram_n_273, B1 => gl_ram_n_430, B2 => gl_ram_ram_31(1), C => n_0, Z => gl_ram_n_572);
  gl_ram_g28308 : AO221D0BWP7T port map(A1 => gl_ram_n_476, A2 => gl_ram_n_277, B1 => gl_ram_n_414, B2 => gl_ram_ram_0(0), C => n_0, Z => gl_ram_n_571);
  gl_ram_g28309 : AO221D0BWP7T port map(A1 => gl_ram_n_491, A2 => gl_ram_n_273, B1 => gl_ram_n_430, B2 => gl_ram_ram_31(2), C => n_0, Z => gl_ram_n_570);
  gl_ram_g28310 : AO221D0BWP7T port map(A1 => gl_ram_n_476, A2 => gl_ram_n_281, B1 => gl_ram_n_435, B2 => gl_ram_ram_32(0), C => n_0, Z => gl_ram_n_569);
  gl_ram_g28311 : AO221D0BWP7T port map(A1 => gl_ram_n_488, A2 => gl_ram_n_281, B1 => gl_ram_n_435, B2 => gl_ram_ram_32(1), C => n_0, Z => gl_ram_n_568);
  gl_ram_g28312 : AO221D0BWP7T port map(A1 => gl_ram_n_475, A2 => gl_ram_n_281, B1 => gl_ram_n_435, B2 => gl_ram_ram_32(2), C => n_0, Z => gl_ram_n_567);
  gl_ram_g28313 : AO221D0BWP7T port map(A1 => gl_ram_n_476, A2 => gl_ram_n_283, B1 => gl_ram_n_387, B2 => gl_ram_ram_33(0), C => n_0, Z => gl_ram_n_566);
  gl_ram_g28314 : AO221D0BWP7T port map(A1 => gl_ram_n_488, A2 => gl_ram_n_283, B1 => gl_ram_n_387, B2 => gl_ram_ram_33(1), C => n_0, Z => gl_ram_n_565);
  gl_ram_g28315 : AO221D0BWP7T port map(A1 => gl_ram_n_475, A2 => gl_ram_n_283, B1 => gl_ram_n_387, B2 => gl_ram_ram_33(2), C => n_0, Z => gl_ram_n_564);
  gl_ram_g28316 : AO221D0BWP7T port map(A1 => gl_ram_n_476, A2 => gl_ram_n_280, B1 => gl_ram_n_419, B2 => gl_ram_ram_34(0), C => n_0, Z => gl_ram_n_563);
  gl_ram_g28317 : AO221D0BWP7T port map(A1 => gl_ram_n_488, A2 => gl_ram_n_280, B1 => gl_ram_n_419, B2 => gl_ram_ram_34(1), C => n_0, Z => gl_ram_n_562);
  gl_ram_g28318 : AO221D0BWP7T port map(A1 => gl_ram_n_475, A2 => gl_ram_n_280, B1 => gl_ram_n_419, B2 => gl_ram_ram_34(2), C => n_0, Z => gl_ram_n_561);
  gl_ram_g28319 : AO221D0BWP7T port map(A1 => gl_ram_n_476, A2 => gl_ram_n_282, B1 => gl_ram_n_364, B2 => gl_ram_ram_35(0), C => n_0, Z => gl_ram_n_560);
  gl_ram_g28320 : AO221D0BWP7T port map(A1 => gl_ram_n_488, A2 => gl_ram_n_282, B1 => gl_ram_n_364, B2 => gl_ram_ram_35(1), C => n_0, Z => gl_ram_n_559);
  gl_ram_g28321 : AO221D0BWP7T port map(A1 => gl_ram_n_475, A2 => gl_ram_n_282, B1 => gl_ram_n_364, B2 => gl_ram_ram_35(2), C => n_0, Z => gl_ram_n_558);
  gl_ram_g28322 : AO221D0BWP7T port map(A1 => gl_ram_n_478, A2 => gl_ram_n_281, B1 => gl_ram_n_422, B2 => gl_ram_ram_36(0), C => n_0, Z => gl_ram_n_557);
  gl_ram_g28323 : AO221D0BWP7T port map(A1 => gl_ram_n_493, A2 => gl_ram_n_281, B1 => gl_ram_n_422, B2 => gl_ram_ram_36(1), C => n_0, Z => gl_ram_n_556);
  gl_ram_g28324 : AO221D0BWP7T port map(A1 => gl_ram_n_477, A2 => gl_ram_n_281, B1 => gl_ram_n_422, B2 => gl_ram_ram_36(2), C => n_0, Z => gl_ram_n_555);
  gl_ram_g28325 : AO221D0BWP7T port map(A1 => gl_ram_n_478, A2 => gl_ram_n_283, B1 => gl_ram_n_386, B2 => gl_ram_ram_37(0), C => n_0, Z => gl_ram_n_554);
  gl_ram_g28326 : AO221D0BWP7T port map(A1 => gl_ram_n_493, A2 => gl_ram_n_283, B1 => gl_ram_n_386, B2 => gl_ram_ram_37(1), C => n_0, Z => gl_ram_n_553);
  gl_ram_g28327 : AO221D0BWP7T port map(A1 => gl_ram_n_477, A2 => gl_ram_n_283, B1 => gl_ram_n_386, B2 => gl_ram_ram_37(2), C => n_0, Z => gl_ram_n_552);
  gl_ram_g28328 : AO221D0BWP7T port map(A1 => gl_ram_n_478, A2 => gl_ram_n_280, B1 => gl_ram_n_394, B2 => gl_ram_ram_38(0), C => n_0, Z => gl_ram_n_551);
  gl_ram_g28329 : AO221D0BWP7T port map(A1 => gl_ram_n_493, A2 => gl_ram_n_280, B1 => gl_ram_n_394, B2 => gl_ram_ram_38(1), C => n_0, Z => gl_ram_n_550);
  gl_ram_g28330 : AO221D0BWP7T port map(A1 => gl_ram_n_477, A2 => gl_ram_n_280, B1 => gl_ram_n_394, B2 => gl_ram_ram_38(2), C => n_0, Z => gl_ram_n_549);
  gl_ram_g28331 : AO221D0BWP7T port map(A1 => gl_ram_n_475, A2 => gl_ram_n_277, B1 => gl_ram_n_414, B2 => gl_ram_ram_0(2), C => n_0, Z => gl_ram_n_548);
  gl_ram_g28332 : AO221D0BWP7T port map(A1 => gl_ram_n_478, A2 => gl_ram_n_282, B1 => gl_ram_n_379, B2 => gl_ram_ram_39(0), C => n_0, Z => gl_ram_n_547);
  gl_ram_g28333 : AO221D0BWP7T port map(A1 => gl_ram_n_493, A2 => gl_ram_n_282, B1 => gl_ram_n_379, B2 => gl_ram_ram_39(1), C => n_0, Z => gl_ram_n_546);
  gl_ram_g28334 : AO221D0BWP7T port map(A1 => gl_ram_n_477, A2 => gl_ram_n_282, B1 => gl_ram_n_379, B2 => gl_ram_ram_39(2), C => n_0, Z => gl_ram_n_545);
  gl_ram_g28335 : AO221D0BWP7T port map(A1 => gl_ram_n_476, A2 => gl_ram_n_287, B1 => gl_ram_n_441, B2 => gl_ram_ram_40(0), C => n_0, Z => gl_ram_n_544);
  gl_ram_g28336 : AO221D0BWP7T port map(A1 => gl_ram_n_488, A2 => gl_ram_n_287, B1 => gl_ram_n_441, B2 => gl_ram_ram_40(1), C => n_0, Z => gl_ram_n_543);
  gl_ram_g28337 : AO221D0BWP7T port map(A1 => gl_ram_n_475, A2 => gl_ram_n_287, B1 => gl_ram_n_441, B2 => gl_ram_ram_40(2), C => n_0, Z => gl_ram_n_542);
  gl_ram_g28338 : AO221D0BWP7T port map(A1 => gl_ram_n_488, A2 => gl_ram_n_285, B1 => gl_ram_n_401, B2 => gl_ram_ram_41(1), C => n_0, Z => gl_ram_n_541);
  gl_ram_g28339 : AO221D0BWP7T port map(A1 => gl_ram_n_476, A2 => gl_ram_n_285, B1 => gl_ram_n_401, B2 => gl_ram_ram_41(0), C => n_0, Z => gl_ram_n_540);
  gl_ram_g28340 : AO221D0BWP7T port map(A1 => gl_ram_n_475, A2 => gl_ram_n_285, B1 => gl_ram_n_401, B2 => gl_ram_ram_41(2), C => n_0, Z => gl_ram_n_539);
  gl_ram_g28341 : AO221D0BWP7T port map(A1 => gl_ram_n_476, A2 => gl_ram_n_286, B1 => gl_ram_n_389, B2 => gl_ram_ram_42(0), C => n_0, Z => gl_ram_n_538);
  gl_ram_g28342 : AO221D0BWP7T port map(A1 => gl_ram_n_488, A2 => gl_ram_n_286, B1 => gl_ram_n_389, B2 => gl_ram_ram_42(1), C => n_0, Z => gl_ram_n_537);
  gl_ram_g28343 : AO221D0BWP7T port map(A1 => gl_ram_n_476, A2 => gl_ram_n_284, B1 => gl_ram_n_357, B2 => gl_ram_ram_43(0), C => n_0, Z => gl_ram_n_536);
  gl_ram_g28344 : AO221D0BWP7T port map(A1 => gl_ram_n_475, A2 => gl_ram_n_286, B1 => gl_ram_n_389, B2 => gl_ram_ram_42(2), C => n_0, Z => gl_ram_n_535);
  gl_ram_g28345 : AO221D0BWP7T port map(A1 => gl_ram_n_488, A2 => gl_ram_n_284, B1 => gl_ram_n_357, B2 => gl_ram_ram_43(1), C => n_0, Z => gl_ram_n_534);
  gl_ram_g28346 : AO221D0BWP7T port map(A1 => gl_ram_n_475, A2 => gl_ram_n_284, B1 => gl_ram_n_357, B2 => gl_ram_ram_43(2), C => n_0, Z => gl_ram_n_533);
  gl_ram_g28347 : AO221D0BWP7T port map(A1 => gl_ram_n_478, A2 => gl_ram_n_287, B1 => gl_ram_n_429, B2 => gl_ram_ram_44(0), C => n_0, Z => gl_ram_n_532);
  gl_ram_g28348 : AO221D0BWP7T port map(A1 => gl_ram_n_493, A2 => gl_ram_n_287, B1 => gl_ram_n_429, B2 => gl_ram_ram_44(1), C => n_0, Z => gl_ram_n_531);
  gl_ram_g28349 : AO221D0BWP7T port map(A1 => gl_ram_n_477, A2 => gl_ram_n_287, B1 => gl_ram_n_429, B2 => gl_ram_ram_44(2), C => n_0, Z => gl_ram_n_530);
  gl_ram_g28350 : AO221D0BWP7T port map(A1 => gl_ram_n_478, A2 => gl_ram_n_285, B1 => gl_ram_n_399, B2 => gl_ram_ram_45(0), C => n_0, Z => gl_ram_n_529);
  gl_ram_g28351 : AO221D0BWP7T port map(A1 => gl_ram_n_493, A2 => gl_ram_n_285, B1 => gl_ram_n_399, B2 => gl_ram_ram_45(1), C => n_0, Z => gl_ram_n_528);
  gl_ram_g28352 : AO221D0BWP7T port map(A1 => gl_ram_n_477, A2 => gl_ram_n_285, B1 => gl_ram_n_399, B2 => gl_ram_ram_45(2), C => n_0, Z => gl_ram_n_527);
  gl_ram_g28353 : AO221D0BWP7T port map(A1 => gl_ram_n_478, A2 => gl_ram_n_286, B1 => gl_ram_n_396, B2 => gl_ram_ram_46(0), C => n_0, Z => gl_ram_n_526);
  gl_ram_g28354 : AO221D0BWP7T port map(A1 => gl_ram_n_493, A2 => gl_ram_n_286, B1 => gl_ram_n_396, B2 => gl_ram_ram_46(1), C => n_0, Z => gl_ram_n_525);
  gl_ram_g28355 : AO221D0BWP7T port map(A1 => gl_ram_n_477, A2 => gl_ram_n_286, B1 => gl_ram_n_396, B2 => gl_ram_ram_46(2), C => n_0, Z => gl_ram_n_524);
  gl_ram_g28356 : AO221D0BWP7T port map(A1 => gl_ram_n_478, A2 => gl_ram_n_284, B1 => gl_ram_n_378, B2 => gl_ram_ram_47(0), C => n_0, Z => gl_ram_n_523);
  gl_ram_g28357 : AO221D0BWP7T port map(A1 => gl_ram_n_493, A2 => gl_ram_n_284, B1 => gl_ram_n_378, B2 => gl_ram_ram_47(1), C => n_0, Z => gl_ram_n_522);
  gl_ram_g28358 : AO221D0BWP7T port map(A1 => gl_ram_n_477, A2 => gl_ram_n_284, B1 => gl_ram_n_378, B2 => gl_ram_ram_47(2), C => n_0, Z => gl_ram_n_521);
  gl_ram_g28359 : AO221D0BWP7T port map(A1 => gl_ram_n_473, A2 => gl_ram_n_281, B1 => gl_ram_n_393, B2 => gl_ram_ram_48(0), C => n_0, Z => gl_ram_n_520);
  gl_ram_g28360 : AO221D0BWP7T port map(A1 => gl_ram_n_492, A2 => gl_ram_n_281, B1 => gl_ram_n_393, B2 => gl_ram_ram_48(1), C => n_0, Z => gl_ram_n_519);
  gl_ram_g28361 : AO221D0BWP7T port map(A1 => gl_ram_n_474, A2 => gl_ram_n_281, B1 => gl_ram_n_393, B2 => gl_ram_ram_48(2), C => n_0, Z => gl_ram_n_518);
  gl_ram_g28362 : AO221D0BWP7T port map(A1 => gl_ram_n_473, A2 => gl_ram_n_283, B1 => gl_ram_n_398, B2 => gl_ram_ram_49(0), C => n_0, Z => gl_ram_n_517);
  gl_ram_g28363 : AO221D0BWP7T port map(A1 => gl_ram_n_492, A2 => gl_ram_n_283, B1 => gl_ram_n_398, B2 => gl_ram_ram_49(1), C => n_0, Z => gl_ram_n_516);
  gl_ram_g28364 : AO221D0BWP7T port map(A1 => gl_ram_n_474, A2 => gl_ram_n_283, B1 => gl_ram_n_398, B2 => gl_ram_ram_49(2), C => n_0, Z => gl_ram_n_515);
  gl_ram_g28365 : AO221D0BWP7T port map(A1 => gl_ram_n_473, A2 => gl_ram_n_280, B1 => gl_ram_n_367, B2 => gl_ram_ram_50(0), C => n_0, Z => gl_ram_n_514);
  gl_ram_g28366 : AO221D0BWP7T port map(A1 => gl_ram_n_492, A2 => gl_ram_n_280, B1 => gl_ram_n_367, B2 => gl_ram_ram_50(1), C => n_0, Z => gl_ram_n_513);
  gl_ram_g28367 : AO221D0BWP7T port map(A1 => gl_ram_n_474, A2 => gl_ram_n_280, B1 => gl_ram_n_367, B2 => gl_ram_ram_50(2), C => n_0, Z => gl_ram_n_512);
  gl_ram_g28368 : AO221D0BWP7T port map(A1 => gl_ram_n_473, A2 => gl_ram_n_282, B1 => gl_ram_n_397, B2 => gl_ram_ram_51(0), C => n_0, Z => gl_ram_n_511);
  gl_ram_g28369 : AO221D0BWP7T port map(A1 => gl_ram_n_492, A2 => gl_ram_n_282, B1 => gl_ram_n_397, B2 => gl_ram_ram_51(1), C => n_0, Z => gl_ram_n_510);
  gl_ram_g28370 : AO221D0BWP7T port map(A1 => gl_ram_n_474, A2 => gl_ram_n_282, B1 => gl_ram_n_397, B2 => gl_ram_ram_51(2), C => n_0, Z => gl_ram_n_509);
  gl_ram_g28371 : AO221D0BWP7T port map(A1 => gl_ram_n_489, A2 => gl_ram_n_281, B1 => gl_ram_n_385, B2 => gl_ram_ram_52(0), C => n_0, Z => gl_ram_n_508);
  gl_ram_g28372 : AO221D0BWP7T port map(A1 => gl_ram_n_490, A2 => gl_ram_n_281, B1 => gl_ram_n_385, B2 => gl_ram_ram_52(1), C => n_0, Z => gl_ram_n_507);
  gl_ram_g28373 : AO221D0BWP7T port map(A1 => gl_ram_n_491, A2 => gl_ram_n_281, B1 => gl_ram_n_385, B2 => gl_ram_ram_52(2), C => n_0, Z => gl_ram_n_506);
  gl_ram_g28374 : AO221D0BWP7T port map(A1 => gl_ram_n_489, A2 => gl_ram_n_283, B1 => gl_ram_n_369, B2 => gl_ram_ram_53(0), C => n_0, Z => gl_ram_n_505);
  gl_ram_g28375 : AO221D0BWP7T port map(A1 => gl_ram_n_490, A2 => gl_ram_n_283, B1 => gl_ram_n_369, B2 => gl_ram_ram_53(1), C => n_0, Z => gl_ram_n_504);
  gl_ram_g28376 : AO221D0BWP7T port map(A1 => gl_ram_n_491, A2 => gl_ram_n_283, B1 => gl_ram_n_369, B2 => gl_ram_ram_53(2), C => n_0, Z => gl_ram_n_503);
  gl_ram_g28377 : AO221D0BWP7T port map(A1 => gl_ram_n_489, A2 => gl_ram_n_280, B1 => gl_ram_n_363, B2 => gl_ram_ram_54(0), C => n_0, Z => gl_ram_n_502);
  gl_ram_g28378 : AO221D0BWP7T port map(A1 => gl_ram_n_490, A2 => gl_ram_n_280, B1 => gl_ram_n_363, B2 => gl_ram_ram_54(1), C => n_0, Z => gl_ram_n_501);
  gl_ram_g28379 : AO22D0BWP7T port map(A1 => gl_ram_n_487, A2 => gl_ram_n_324, B1 => gl_ram_ram_position(5), B2 => gl_ram_n_0, Z => gl_ram_n_500);
  gl_ram_g28380 : XNR2D1BWP7T port map(A1 => gl_ram_n_486, A2 => gl_ram_y_grid(3), ZN => gl_ram_n_499);
  gl_ram_g28381 : FA1D0BWP7T port map(A => gl_ram_n_56, B => gl_ram_y_grid(2), CI => gl_ram_n_466, CO => gl_ram_n_486, S => gl_ram_n_487);
  gl_ram_g28382 : NR2D1BWP7T port map(A1 => gl_ram_n_471, A2 => gl_ram_n_350, ZN => gl_ram_n_498);
  gl_ram_g28383 : NR2D1BWP7T port map(A1 => gl_ram_n_471, A2 => gl_ram_n_343, ZN => gl_ram_n_497);
  gl_ram_g28384 : AN2D1BWP7T port map(A1 => gl_ram_n_472, A2 => gl_ram_n_344, Z => gl_ram_n_496);
  gl_ram_g28385 : NR2D1BWP7T port map(A1 => gl_ram_n_470, A2 => gl_ram_n_345, ZN => gl_ram_n_495);
  gl_ram_g28386 : NR2D1BWP7T port map(A1 => gl_ram_n_469, A2 => gl_ram_n_345, ZN => gl_ram_n_494);
  gl_ram_g28387 : AN2D1BWP7T port map(A1 => gl_ram_n_472, A2 => gl_ram_n_349, Z => gl_ram_n_493);
  gl_ram_g28388 : AN2D1BWP7T port map(A1 => gl_ram_n_472, A2 => gl_ram_n_348, Z => gl_ram_n_492);
  gl_ram_g28389 : NR2XD0BWP7T port map(A1 => gl_ram_n_469, A2 => gl_ram_n_347, ZN => gl_ram_n_491);
  gl_ram_g28390 : AN2D1BWP7T port map(A1 => gl_ram_n_472, A2 => gl_ram_n_346, Z => gl_ram_n_490);
  gl_ram_g28391 : NR2XD0BWP7T port map(A1 => gl_ram_n_470, A2 => gl_ram_n_347, ZN => gl_ram_n_489);
  gl_ram_g28392 : NR2XD0BWP7T port map(A1 => gl_ram_n_471, A2 => gl_ram_n_342, ZN => gl_ram_n_488);
  gl_ram_g28394 : NR2D1BWP7T port map(A1 => gl_ram_n_470, A2 => gl_ram_n_350, ZN => gl_ram_n_485);
  gl_ram_g28395 : NR2D1BWP7T port map(A1 => gl_ram_n_469, A2 => gl_ram_n_350, ZN => gl_ram_n_484);
  gl_ram_g28396 : NR2D1BWP7T port map(A1 => gl_ram_n_469, A2 => gl_ram_n_343, ZN => gl_ram_n_483);
  gl_ram_g28397 : NR2D1BWP7T port map(A1 => gl_ram_n_470, A2 => gl_ram_n_343, ZN => gl_ram_n_482);
  gl_ram_g28398 : NR2XD0BWP7T port map(A1 => gl_ram_n_469, A2 => gl_ram_n_341, ZN => gl_ram_n_481);
  gl_ram_g28399 : NR2XD0BWP7T port map(A1 => gl_ram_n_471, A2 => gl_ram_n_341, ZN => gl_ram_n_480);
  gl_ram_g28400 : NR2XD0BWP7T port map(A1 => gl_ram_n_470, A2 => gl_ram_n_341, ZN => gl_ram_n_479);
  gl_ram_g28401 : INR2XD0BWP7T port map(A1 => gl_ram_n_349, B1 => gl_ram_n_470, ZN => gl_ram_n_478);
  gl_ram_g28402 : INR2XD0BWP7T port map(A1 => gl_ram_n_349, B1 => gl_ram_n_469, ZN => gl_ram_n_477);
  gl_ram_g28403 : NR2XD0BWP7T port map(A1 => gl_ram_n_470, A2 => gl_ram_n_342, ZN => gl_ram_n_476);
  gl_ram_g28404 : NR2XD0BWP7T port map(A1 => gl_ram_n_469, A2 => gl_ram_n_342, ZN => gl_ram_n_475);
  gl_ram_g28405 : INR2XD0BWP7T port map(A1 => gl_ram_n_348, B1 => gl_ram_n_469, ZN => gl_ram_n_474);
  gl_ram_g28406 : INR2XD0BWP7T port map(A1 => gl_ram_n_348, B1 => gl_ram_n_470, ZN => gl_ram_n_473);
  gl_ram_g28407 : INVD1BWP7T port map(I => gl_ram_n_472, ZN => gl_ram_n_471);
  gl_ram_g28408 : OAI211D1BWP7T port map(A1 => gl_ram_n_50, A2 => gl_ram_n_319, B => gl_ram_n_462, C => gl_ram_n_6, ZN => gl_ram_n_472);
  gl_ram_g28409 : AOI211XD0BWP7T port map(A1 => gl_ram_n_318, A2 => gl_ram_n_35, B => gl_ram_n_464, C => sig_middelsteknop, ZN => gl_ram_n_470);
  gl_ram_g28410 : AO22D0BWP7T port map(A1 => gl_ram_n_467, A2 => gl_ram_n_324, B1 => gl_ram_ram_position(4), B2 => gl_ram_n_0, Z => gl_ram_n_468);
  gl_ram_g28411 : AOI211XD0BWP7T port map(A1 => gl_ram_n_317, A2 => gl_ram_n_35, B => gl_ram_n_463, C => sig_middelsteknop, ZN => gl_ram_n_469);
  gl_ram_g28424 : FA1D0BWP7T port map(A => gl_ram_n_57, B => gl_ram_n_54, CI => gl_ram_n_312, CO => gl_ram_n_466, S => gl_ram_n_467);
  gl_ram_g28425 : AO22D0BWP7T port map(A1 => gl_ram_n_313, A2 => gl_ram_n_324, B1 => gl_ram_ram_position(3), B2 => gl_ram_n_0, Z => gl_ram_n_465);
  gl_ram_g28426 : MOAI22D0BWP7T port map(A1 => gl_ram_n_320, A2 => gl_ram_n_50, B1 => sig_output_color(0), B2 => gl_ram_n_7, ZN => gl_ram_n_464);
  gl_ram_g28427 : MOAI22D0BWP7T port map(A1 => gl_ram_n_321, A2 => gl_ram_n_50, B1 => sig_output_color(2), B2 => gl_ram_n_7, ZN => gl_ram_n_463);
  gl_ram_g28428 : AOI22D0BWP7T port map(A1 => gl_ram_n_322, A2 => gl_ram_n_35, B1 => sig_output_color(1), B2 => gl_ram_n_7, ZN => gl_ram_n_462);
  gl_ram_g28429 : AO22D0BWP7T port map(A1 => gl_ram_n_324, A2 => sig_logic_y(0), B1 => gl_ram_y_grid(0), B2 => gl_ram_n_0, Z => gl_ram_n_461);
  gl_ram_g28430 : AO22D0BWP7T port map(A1 => gl_ram_n_324, A2 => sig_logic_y(1), B1 => gl_ram_y_grid(1), B2 => gl_ram_n_0, Z => gl_ram_n_460);
  gl_ram_g28431 : AO32D1BWP7T port map(A1 => gl_ram_n_324, A2 => gl_ram_n_209, A3 => sig_logic_x(3), B1 => gl_ram_n_0, B2 => gl_ram_x_grid(3), Z => gl_ram_n_459);
  gl_ram_g28432 : MOAI22D0BWP7T port map(A1 => gl_ram_n_323, A2 => gl_ram_n_26, B1 => gl_ram_n_0, B2 => gl_ram_x_grid(1), ZN => gl_ram_n_458);
  gl_ram_g28433 : AO22D0BWP7T port map(A1 => gl_ram_n_324, A2 => gl_ram_x_grid(0), B1 => gl_ram_ram_position(0), B2 => gl_ram_n_0, Z => gl_ram_n_457);
  gl_ram_g28434 : MOAI22D0BWP7T port map(A1 => gl_ram_n_323, A2 => gl_ram_n_220, B1 => gl_ram_n_0, B2 => gl_ram_x_grid(2), ZN => gl_ram_n_456);
  gl_ram_g28435 : MOAI22D0BWP7T port map(A1 => gl_ram_n_323, A2 => gl_ram_n_27, B1 => gl_ram_n_0, B2 => gl_ram_ram_position(1), ZN => gl_ram_n_455);
  gl_ram_g28436 : AO22D0BWP7T port map(A1 => gl_ram_n_324, A2 => gl_ram_n_271, B1 => gl_ram_ram_position(2), B2 => gl_ram_n_0, Z => gl_ram_n_454);
  gl_ram_g28437 : MOAI22D0BWP7T port map(A1 => gl_ram_n_323, A2 => sig_logic_x(0), B1 => gl_ram_n_0, B2 => gl_ram_x_grid(0), ZN => gl_ram_n_453);
  gl_ram_g28438 : MOAI22D0BWP7T port map(A1 => gl_ram_n_323, A2 => sig_logic_y(2), B1 => gl_ram_n_0, B2 => gl_ram_y_grid(2), ZN => gl_ram_n_452);
  gl_ram_g28439 : MOAI22D0BWP7T port map(A1 => gl_ram_n_323, A2 => gl_ram_n_22, B1 => gl_ram_n_0, B2 => gl_ram_y_grid(3), ZN => gl_ram_n_451);
  gl_ram_g28440 : ND2D1BWP7T port map(A1 => gl_ram_n_223, A2 => gl_ram_n_338, ZN => gl_ram_n_450);
  gl_ram_g28441 : ND2D1BWP7T port map(A1 => gl_ram_n_223, A2 => gl_ram_n_337, ZN => gl_ram_n_449);
  gl_ram_g28442 : ND2D1BWP7T port map(A1 => gl_ram_n_222, A2 => gl_ram_n_337, ZN => gl_ram_n_448);
  gl_ram_g28443 : ND2D1BWP7T port map(A1 => gl_ram_n_225, A2 => gl_ram_n_337, ZN => gl_ram_n_447);
  gl_ram_g28444 : ND2D1BWP7T port map(A1 => gl_ram_n_226, A2 => gl_ram_n_339, ZN => gl_ram_n_446);
  gl_ram_g28445 : ND2D1BWP7T port map(A1 => gl_ram_n_225, A2 => gl_ram_n_339, ZN => gl_ram_n_445);
  gl_ram_g28446 : ND2D1BWP7T port map(A1 => gl_ram_n_223, A2 => gl_ram_n_340, ZN => gl_ram_n_444);
  gl_ram_g28447 : ND2D1BWP7T port map(A1 => gl_ram_n_227, A2 => gl_ram_n_335, ZN => gl_ram_n_443);
  gl_ram_g28448 : ND2D1BWP7T port map(A1 => gl_ram_n_226, A2 => gl_ram_n_338, ZN => gl_ram_n_442);
  gl_ram_g28449 : ND2D1BWP7T port map(A1 => gl_ram_n_334, A2 => gl_ram_n_229, ZN => gl_ram_n_441);
  gl_ram_g28450 : ND2D1BWP7T port map(A1 => gl_ram_n_225, A2 => gl_ram_n_340, ZN => gl_ram_n_440);
  gl_ram_g28451 : ND2D1BWP7T port map(A1 => gl_ram_n_226, A2 => gl_ram_n_340, ZN => gl_ram_n_439);
  gl_ram_g28452 : ND2D1BWP7T port map(A1 => gl_ram_n_223, A2 => gl_ram_n_339, ZN => gl_ram_n_438);
  gl_ram_g28453 : ND2D1BWP7T port map(A1 => gl_ram_n_222, A2 => gl_ram_n_340, ZN => gl_ram_n_437);
  gl_ram_g28454 : ND2D1BWP7T port map(A1 => gl_ram_n_222, A2 => gl_ram_n_339, ZN => gl_ram_n_436);
  gl_ram_g28455 : ND2D1BWP7T port map(A1 => gl_ram_n_334, A2 => gl_ram_n_227, ZN => gl_ram_n_435);
  gl_ram_g28456 : ND2D1BWP7T port map(A1 => gl_ram_n_225, A2 => gl_ram_n_338, ZN => gl_ram_n_434);
  gl_ram_g28457 : ND2D1BWP7T port map(A1 => gl_ram_n_223, A2 => gl_ram_n_336, ZN => gl_ram_n_433);
  gl_ram_g28458 : ND2D1BWP7T port map(A1 => gl_ram_n_228, A2 => gl_ram_n_335, ZN => gl_ram_n_432);
  gl_ram_g28459 : ND2D1BWP7T port map(A1 => gl_ram_n_226, A2 => gl_ram_n_331, ZN => gl_ram_n_431);
  gl_ram_g28460 : ND2D1BWP7T port map(A1 => gl_ram_n_226, A2 => gl_ram_n_330, ZN => gl_ram_n_430);
  gl_ram_g28461 : ND2D1BWP7T port map(A1 => gl_ram_n_333, A2 => gl_ram_n_229, ZN => gl_ram_n_429);
  gl_ram_g28462 : ND2D1BWP7T port map(A1 => gl_ram_n_223, A2 => gl_ram_n_335, ZN => gl_ram_n_428);
  gl_ram_g28463 : ND2D1BWP7T port map(A1 => gl_ram_n_225, A2 => gl_ram_n_336, ZN => gl_ram_n_427);
  gl_ram_g28464 : ND2D1BWP7T port map(A1 => gl_ram_n_222, A2 => gl_ram_n_338, ZN => gl_ram_n_426);
  gl_ram_g28465 : ND2D1BWP7T port map(A1 => gl_ram_n_226, A2 => gl_ram_n_336, ZN => gl_ram_n_425);
  gl_ram_g28466 : ND2D1BWP7T port map(A1 => gl_ram_n_222, A2 => gl_ram_n_336, ZN => gl_ram_n_424);
  gl_ram_g28467 : ND2D1BWP7T port map(A1 => gl_ram_n_226, A2 => gl_ram_n_337, ZN => gl_ram_n_423);
  gl_ram_g28468 : ND2D1BWP7T port map(A1 => gl_ram_n_333, A2 => gl_ram_n_227, ZN => gl_ram_n_422);
  gl_ram_g28469 : ND2D1BWP7T port map(A1 => gl_ram_n_225, A2 => gl_ram_n_331, ZN => gl_ram_n_421);
  gl_ram_g28470 : ND2D1BWP7T port map(A1 => gl_ram_n_225, A2 => gl_ram_n_330, ZN => gl_ram_n_420);
  gl_ram_g28471 : ND2D1BWP7T port map(A1 => gl_ram_n_334, A2 => gl_ram_n_228, ZN => gl_ram_n_419);
  gl_ram_g28472 : ND2D1BWP7T port map(A1 => gl_ram_n_225, A2 => gl_ram_n_335, ZN => gl_ram_n_418);
  gl_ram_g28473 : ND2D1BWP7T port map(A1 => gl_ram_n_226, A2 => gl_ram_n_335, ZN => gl_ram_n_417);
  gl_ram_g28474 : ND2D1BWP7T port map(A1 => gl_ram_n_222, A2 => gl_ram_n_335, ZN => gl_ram_n_416);
  gl_ram_g28475 : ND2D1BWP7T port map(A1 => gl_ram_n_226, A2 => gl_ram_n_332, ZN => gl_ram_n_415);
  gl_ram_g28476 : ND2D1BWP7T port map(A1 => gl_ram_n_223, A2 => gl_ram_n_334, ZN => gl_ram_n_414);
  gl_ram_g28477 : ND2D1BWP7T port map(A1 => gl_ram_n_327, A2 => gl_ram_n_229, ZN => gl_ram_n_413);
  gl_ram_g28478 : ND2D1BWP7T port map(A1 => gl_ram_n_227, A2 => gl_ram_n_328, ZN => gl_ram_n_412);
  gl_ram_g28479 : ND2D1BWP7T port map(A1 => gl_ram_n_226, A2 => gl_ram_n_329, ZN => gl_ram_n_411);
  gl_ram_g28480 : ND2D1BWP7T port map(A1 => gl_ram_n_330, A2 => gl_ram_n_228, ZN => gl_ram_n_410);
  gl_ram_g28481 : ND2D1BWP7T port map(A1 => gl_ram_n_331, A2 => gl_ram_n_229, ZN => gl_ram_n_409);
  gl_ram_g28482 : ND2D1BWP7T port map(A1 => gl_ram_n_331, A2 => gl_ram_n_224, ZN => gl_ram_n_408);
  gl_ram_g28483 : ND2D1BWP7T port map(A1 => gl_ram_n_325, A2 => gl_ram_n_229, ZN => gl_ram_n_407);
  gl_ram_g28484 : ND2D1BWP7T port map(A1 => gl_ram_n_330, A2 => gl_ram_n_224, ZN => gl_ram_n_406);
  gl_ram_g28485 : ND2D1BWP7T port map(A1 => gl_ram_n_330, A2 => gl_ram_n_229, ZN => gl_ram_n_405);
  gl_ram_g28486 : ND2D1BWP7T port map(A1 => gl_ram_n_223, A2 => gl_ram_n_331, ZN => gl_ram_n_404);
  gl_ram_g28487 : ND2D1BWP7T port map(A1 => gl_ram_n_223, A2 => gl_ram_n_330, ZN => gl_ram_n_403);
  gl_ram_g28488 : ND2D1BWP7T port map(A1 => gl_ram_n_222, A2 => gl_ram_n_331, ZN => gl_ram_n_402);
  gl_ram_g28489 : ND2D1BWP7T port map(A1 => gl_ram_n_326, A2 => gl_ram_n_229, ZN => gl_ram_n_401);
  gl_ram_g28490 : ND2D1BWP7T port map(A1 => gl_ram_n_222, A2 => gl_ram_n_330, ZN => gl_ram_n_400);
  gl_ram_g28491 : ND2D1BWP7T port map(A1 => gl_ram_n_332, A2 => gl_ram_n_229, ZN => gl_ram_n_399);
  gl_ram_g28492 : ND2D1BWP7T port map(A1 => gl_ram_n_331, A2 => gl_ram_n_227, ZN => gl_ram_n_398);
  gl_ram_g28493 : ND2D1BWP7T port map(A1 => gl_ram_n_331, A2 => gl_ram_n_228, ZN => gl_ram_n_397);
  gl_ram_g28494 : INVD1BWP7T port map(I => gl_ram_n_346, ZN => gl_ram_n_347);
  gl_ram_g28495 : INVD1BWP7T port map(I => gl_ram_n_344, ZN => gl_ram_n_345);
  gl_ram_g28496 : ND2D1BWP7T port map(A1 => gl_ram_n_333, A2 => gl_ram_n_224, ZN => gl_ram_n_396);
  gl_ram_g28497 : ND2D1BWP7T port map(A1 => gl_ram_n_225, A2 => gl_ram_n_332, ZN => gl_ram_n_395);
  gl_ram_g28498 : ND2D1BWP7T port map(A1 => gl_ram_n_333, A2 => gl_ram_n_228, ZN => gl_ram_n_394);
  gl_ram_g28499 : ND2D1BWP7T port map(A1 => gl_ram_n_327, A2 => gl_ram_n_227, ZN => gl_ram_n_393);
  gl_ram_g28500 : ND2D1BWP7T port map(A1 => gl_ram_n_222, A2 => gl_ram_n_334, ZN => gl_ram_n_392);
  gl_ram_g28501 : ND2D1BWP7T port map(A1 => gl_ram_n_226, A2 => gl_ram_n_334, ZN => gl_ram_n_391);
  gl_ram_g28502 : ND2D1BWP7T port map(A1 => gl_ram_n_225, A2 => gl_ram_n_334, ZN => gl_ram_n_390);
  gl_ram_g28503 : ND2D1BWP7T port map(A1 => gl_ram_n_334, A2 => gl_ram_n_224, ZN => gl_ram_n_389);
  gl_ram_g28504 : ND2D1BWP7T port map(A1 => gl_ram_n_226, A2 => gl_ram_n_326, ZN => gl_ram_n_388);
  gl_ram_g28505 : ND2D1BWP7T port map(A1 => gl_ram_n_326, A2 => gl_ram_n_227, ZN => gl_ram_n_387);
  gl_ram_g28506 : ND2D1BWP7T port map(A1 => gl_ram_n_332, A2 => gl_ram_n_227, ZN => gl_ram_n_386);
  gl_ram_g28507 : ND2D1BWP7T port map(A1 => gl_ram_n_325, A2 => gl_ram_n_227, ZN => gl_ram_n_385);
  gl_ram_g28508 : ND2D1BWP7T port map(A1 => gl_ram_n_226, A2 => gl_ram_n_325, ZN => gl_ram_n_384);
  gl_ram_g28509 : ND2D1BWP7T port map(A1 => gl_ram_n_223, A2 => gl_ram_n_333, ZN => gl_ram_n_383);
  gl_ram_g28510 : ND2D1BWP7T port map(A1 => gl_ram_n_225, A2 => gl_ram_n_329, ZN => gl_ram_n_382);
  gl_ram_g28511 : ND2D1BWP7T port map(A1 => gl_ram_n_223, A2 => gl_ram_n_332, ZN => gl_ram_n_381);
  gl_ram_g28512 : ND2D1BWP7T port map(A1 => gl_ram_n_222, A2 => gl_ram_n_332, ZN => gl_ram_n_380);
  gl_ram_g28513 : ND2D1BWP7T port map(A1 => gl_ram_n_332, A2 => gl_ram_n_228, ZN => gl_ram_n_379);
  gl_ram_g28514 : ND2D1BWP7T port map(A1 => gl_ram_n_332, A2 => gl_ram_n_224, ZN => gl_ram_n_378);
  gl_ram_g28515 : ND2D1BWP7T port map(A1 => gl_ram_n_225, A2 => gl_ram_n_326, ZN => gl_ram_n_377);
  gl_ram_g28516 : ND2D1BWP7T port map(A1 => gl_ram_n_225, A2 => gl_ram_n_325, ZN => gl_ram_n_376);
  gl_ram_g28517 : ND2D1BWP7T port map(A1 => gl_ram_n_226, A2 => gl_ram_n_328, ZN => gl_ram_n_375);
  gl_ram_g28518 : ND2D1BWP7T port map(A1 => gl_ram_n_226, A2 => gl_ram_n_333, ZN => gl_ram_n_374);
  gl_ram_g28519 : ND2D1BWP7T port map(A1 => gl_ram_n_226, A2 => gl_ram_n_327, ZN => gl_ram_n_373);
  gl_ram_g28520 : ND2D1BWP7T port map(A1 => gl_ram_n_228, A2 => gl_ram_n_328, ZN => gl_ram_n_372);
  gl_ram_g28521 : ND2D1BWP7T port map(A1 => gl_ram_n_225, A2 => gl_ram_n_333, ZN => gl_ram_n_371);
  gl_ram_g28522 : ND2D1BWP7T port map(A1 => gl_ram_n_222, A2 => gl_ram_n_333, ZN => gl_ram_n_370);
  gl_ram_g28523 : ND2D1BWP7T port map(A1 => gl_ram_n_330, A2 => gl_ram_n_227, ZN => gl_ram_n_369);
  gl_ram_g28524 : ND2D1BWP7T port map(A1 => gl_ram_n_223, A2 => gl_ram_n_328, ZN => gl_ram_n_368);
  gl_ram_g28525 : ND2D1BWP7T port map(A1 => gl_ram_n_327, A2 => gl_ram_n_228, ZN => gl_ram_n_367);
  gl_ram_g28526 : ND2D1BWP7T port map(A1 => gl_ram_n_223, A2 => gl_ram_n_329, ZN => gl_ram_n_366);
  gl_ram_g28527 : ND2D1BWP7T port map(A1 => gl_ram_n_222, A2 => gl_ram_n_329, ZN => gl_ram_n_365);
  gl_ram_g28528 : ND2D1BWP7T port map(A1 => gl_ram_n_326, A2 => gl_ram_n_228, ZN => gl_ram_n_364);
  gl_ram_g28529 : ND2D1BWP7T port map(A1 => gl_ram_n_325, A2 => gl_ram_n_228, ZN => gl_ram_n_363);
  gl_ram_g28530 : ND2D1BWP7T port map(A1 => gl_ram_n_223, A2 => gl_ram_n_327, ZN => gl_ram_n_362);
  gl_ram_g28531 : ND2D1BWP7T port map(A1 => gl_ram_n_225, A2 => gl_ram_n_328, ZN => gl_ram_n_361);
  gl_ram_g28532 : ND2D1BWP7T port map(A1 => gl_ram_n_225, A2 => gl_ram_n_327, ZN => gl_ram_n_360);
  gl_ram_g28533 : ND2D1BWP7T port map(A1 => gl_ram_n_223, A2 => gl_ram_n_326, ZN => gl_ram_n_359);
  gl_ram_g28534 : ND2D1BWP7T port map(A1 => gl_ram_n_222, A2 => gl_ram_n_326, ZN => gl_ram_n_358);
  gl_ram_g28535 : ND2D1BWP7T port map(A1 => gl_ram_n_326, A2 => gl_ram_n_224, ZN => gl_ram_n_357);
  gl_ram_g28536 : ND2D1BWP7T port map(A1 => gl_ram_n_325, A2 => gl_ram_n_224, ZN => gl_ram_n_356);
  gl_ram_g28537 : ND2D1BWP7T port map(A1 => gl_ram_n_223, A2 => gl_ram_n_325, ZN => gl_ram_n_355);
  gl_ram_g28538 : ND2D1BWP7T port map(A1 => gl_ram_n_222, A2 => gl_ram_n_325, ZN => gl_ram_n_354);
  gl_ram_g28539 : ND2D1BWP7T port map(A1 => gl_ram_n_222, A2 => gl_ram_n_328, ZN => gl_ram_n_353);
  gl_ram_g28540 : ND2D1BWP7T port map(A1 => gl_ram_n_327, A2 => gl_ram_n_224, ZN => gl_ram_n_352);
  gl_ram_g28541 : ND2D1BWP7T port map(A1 => gl_ram_n_222, A2 => gl_ram_n_327, ZN => gl_ram_n_351);
  gl_ram_g28542 : OAI21D0BWP7T port map(A1 => gl_ram_n_311, A2 => sig_middelsteknop, B => gl_ram_n_17, ZN => gl_ram_n_350);
  gl_ram_g28543 : OAI21D0BWP7T port map(A1 => gl_ram_n_316, A2 => gl_ram_ram_position(4), B => gl_ram_n_6, ZN => gl_ram_n_349);
  gl_ram_g28544 : AOI21D0BWP7T port map(A1 => gl_ram_n_315, A2 => gl_ram_n_6, B => gl_ram_n_18, ZN => gl_ram_n_348);
  gl_ram_g28545 : AOI21D0BWP7T port map(A1 => gl_ram_n_316, A2 => gl_ram_n_6, B => gl_ram_n_18, ZN => gl_ram_n_346);
  gl_ram_g28546 : AOI21D0BWP7T port map(A1 => gl_ram_n_309, A2 => gl_ram_n_6, B => gl_ram_n_18, ZN => gl_ram_n_344);
  gl_ram_g28547 : AOI21D0BWP7T port map(A1 => gl_ram_n_310, A2 => gl_ram_n_1, B => sig_middelsteknop, ZN => gl_ram_n_343);
  gl_ram_g28548 : AOI21D0BWP7T port map(A1 => gl_ram_n_314, A2 => gl_ram_n_1, B => sig_middelsteknop, ZN => gl_ram_n_342);
  gl_ram_g28549 : AOI21D0BWP7T port map(A1 => gl_ram_n_311, A2 => gl_ram_n_1, B => sig_middelsteknop, ZN => gl_ram_n_341);
  gl_ram_g28550 : AN2D1BWP7T port map(A1 => gl_ram_n_310, A2 => gl_ram_n_11, Z => gl_ram_n_340);
  gl_ram_g28551 : INR2XD0BWP7T port map(A1 => gl_ram_n_311, B1 => gl_ram_n_10, ZN => gl_ram_n_339);
  gl_ram_g28552 : NR2XD0BWP7T port map(A1 => gl_ram_n_309, A2 => gl_ram_n_8, ZN => gl_ram_n_338);
  gl_ram_g28553 : NR2XD0BWP7T port map(A1 => gl_ram_n_309, A2 => gl_ram_n_10, ZN => gl_ram_n_337);
  gl_ram_g28554 : CKAN2D1BWP7T port map(A1 => gl_ram_n_311, A2 => gl_ram_n_9, Z => gl_ram_n_336);
  gl_ram_g28555 : CKAN2D1BWP7T port map(A1 => gl_ram_n_311, A2 => gl_ram_n_11, Z => gl_ram_n_335);
  gl_ram_g28556 : CKAN2D1BWP7T port map(A1 => gl_ram_n_314, A2 => gl_ram_n_11, Z => gl_ram_n_334);
  gl_ram_g28557 : INR2XD0BWP7T port map(A1 => gl_ram_n_11, B1 => gl_ram_n_316, ZN => gl_ram_n_333);
  gl_ram_g28558 : NR2XD0BWP7T port map(A1 => gl_ram_n_316, A2 => gl_ram_n_8, ZN => gl_ram_n_332);
  gl_ram_g28559 : NR2XD0BWP7T port map(A1 => gl_ram_n_315, A2 => gl_ram_n_10, ZN => gl_ram_n_331);
  gl_ram_g28560 : NR2XD0BWP7T port map(A1 => gl_ram_n_316, A2 => gl_ram_n_10, ZN => gl_ram_n_330);
  gl_ram_g28561 : INVD1BWP7T port map(I => gl_ram_n_324, ZN => gl_ram_n_323);
  gl_ram_g28562 : ND4D0BWP7T port map(A1 => gl_ram_n_296, A2 => gl_ram_n_295, A3 => gl_ram_n_294, A4 => gl_ram_n_293, ZN => gl_ram_n_322);
  gl_ram_g28563 : AN4D0BWP7T port map(A1 => gl_ram_n_304, A2 => gl_ram_n_292, A3 => gl_ram_n_216, A4 => gl_ram_n_221, Z => gl_ram_n_321);
  gl_ram_g28564 : AN4D0BWP7T port map(A1 => gl_ram_n_289, A2 => gl_ram_n_305, A3 => gl_ram_n_215, A4 => gl_ram_n_217, Z => gl_ram_n_320);
  gl_ram_g28565 : AN4D1BWP7T port map(A1 => gl_ram_n_299, A2 => gl_ram_n_302, A3 => gl_ram_n_218, A4 => gl_ram_n_219, Z => gl_ram_n_319);
  gl_ram_g28566 : ND4D0BWP7T port map(A1 => gl_ram_n_297, A2 => gl_ram_n_301, A3 => gl_ram_n_298, A4 => gl_ram_n_291, ZN => gl_ram_n_318);
  gl_ram_g28567 : ND4D0BWP7T port map(A1 => gl_ram_n_303, A2 => gl_ram_n_290, A3 => gl_ram_n_300, A4 => gl_ram_n_306, ZN => gl_ram_n_317);
  gl_ram_g28568 : CKAN2D1BWP7T port map(A1 => gl_ram_n_310, A2 => gl_ram_n_9, Z => gl_ram_n_329);
  gl_ram_g28569 : INR2XD0BWP7T port map(A1 => gl_ram_n_311, B1 => gl_ram_n_8, ZN => gl_ram_n_328);
  gl_ram_g28570 : CKAN2D1BWP7T port map(A1 => gl_ram_n_314, A2 => gl_ram_n_9, Z => gl_ram_n_327);
  gl_ram_g28571 : NR2XD0BWP7T port map(A1 => gl_ram_n_315, A2 => gl_ram_n_8, ZN => gl_ram_n_326);
  gl_ram_g28572 : INR2XD0BWP7T port map(A1 => gl_ram_n_9, B1 => gl_ram_n_316, ZN => gl_ram_n_325);
  gl_ram_g28573 : NR4D0BWP7T port map(A1 => gl_ram_n_0, A2 => gl_ram_n_288, A3 => gl_ram_n_49, A4 => gl_ram_n_21, ZN => gl_ram_n_324);
  gl_ram_g28574 : INVD0BWP7T port map(I => gl_ram_n_315, ZN => gl_ram_n_314);
  gl_ram_g28575 : FA1D0BWP7T port map(A => gl_ram_n_55, B => gl_ram_y_grid(2), CI => gl_ram_n_270, CO => gl_ram_n_312, S => gl_ram_n_313);
  gl_ram_g28576 : ND2D1BWP7T port map(A1 => gl_ram_n_307, A2 => gl_ram_ram_position(2), ZN => gl_ram_n_316);
  gl_ram_g28577 : CKND2D1BWP7T port map(A1 => gl_ram_n_307, A2 => gl_ram_n_2, ZN => gl_ram_n_315);
  gl_ram_g28578 : INVD1BWP7T port map(I => gl_ram_n_310, ZN => gl_ram_n_309);
  gl_ram_g28579 : NR2XD0BWP7T port map(A1 => gl_ram_n_308, A2 => gl_ram_ram_position(2), ZN => gl_ram_n_311);
  gl_ram_g28580 : NR2XD0BWP7T port map(A1 => gl_ram_n_308, A2 => gl_ram_n_2, ZN => gl_ram_n_310);
  gl_ram_g28581 : AOI22D0BWP7T port map(A1 => gl_ram_n_246, A2 => gl_ram_n_45, B1 => gl_ram_n_260, B2 => gl_ram_n_34, ZN => gl_ram_n_306);
  gl_ram_g28582 : AOI22D0BWP7T port map(A1 => gl_ram_n_261, A2 => gl_ram_n_44, B1 => gl_ram_n_234, B2 => gl_ram_n_45, ZN => gl_ram_n_305);
  gl_ram_g28583 : AOI22D0BWP7T port map(A1 => gl_ram_n_236, A2 => gl_ram_n_44, B1 => gl_ram_n_267, B2 => gl_ram_n_45, ZN => gl_ram_n_304);
  gl_ram_g28584 : AOI22D0BWP7T port map(A1 => gl_ram_n_262, A2 => gl_ram_n_48, B1 => gl_ram_n_268, B2 => gl_ram_n_37, ZN => gl_ram_n_303);
  gl_ram_g28585 : AOI22D0BWP7T port map(A1 => gl_ram_n_250, A2 => gl_ram_n_44, B1 => gl_ram_n_251, B2 => gl_ram_n_45, ZN => gl_ram_n_302);
  gl_ram_g28586 : AOI22D0BWP7T port map(A1 => gl_ram_n_265, A2 => gl_ram_n_37, B1 => gl_ram_n_263, B2 => gl_ram_n_48, ZN => gl_ram_n_301);
  gl_ram_g28587 : AOI22D0BWP7T port map(A1 => gl_ram_n_264, A2 => gl_ram_n_44, B1 => gl_ram_n_241, B2 => gl_ram_n_32, ZN => gl_ram_n_300);
  gl_ram_g28588 : AOI22D0BWP7T port map(A1 => gl_ram_n_253, A2 => gl_ram_n_34, B1 => gl_ram_n_254, B2 => gl_ram_n_33, ZN => gl_ram_n_299);
  gl_ram_g28589 : IND2D1BWP7T port map(A1 => gl_ram_n_288, B1 => gl_ram_ram_position(6), ZN => gl_ram_n_308);
  gl_ram_g28590 : NR2XD0BWP7T port map(A1 => gl_ram_ram_position(6), A2 => gl_ram_n_288, ZN => gl_ram_n_307);
  gl_ram_g28591 : AOI22D0BWP7T port map(A1 => gl_ram_n_256, A2 => gl_ram_n_45, B1 => gl_ram_n_269, B2 => gl_ram_n_34, ZN => gl_ram_n_298);
  gl_ram_g28592 : AOI22D0BWP7T port map(A1 => gl_ram_n_258, A2 => gl_ram_n_33, B1 => gl_ram_n_266, B2 => gl_ram_n_36, ZN => gl_ram_n_297);
  gl_ram_g28593 : AOI22D0BWP7T port map(A1 => gl_ram_n_248, A2 => gl_ram_n_33, B1 => gl_ram_n_249, B2 => gl_ram_n_36, ZN => gl_ram_n_296);
  gl_ram_g28594 : AOI22D0BWP7T port map(A1 => gl_ram_n_259, A2 => gl_ram_n_45, B1 => gl_ram_n_247, B2 => gl_ram_n_34, ZN => gl_ram_n_295);
  gl_ram_g28595 : AOI22D0BWP7T port map(A1 => gl_ram_n_244, A2 => gl_ram_n_37, B1 => gl_ram_n_245, B2 => gl_ram_n_48, ZN => gl_ram_n_294);
  gl_ram_g28596 : AOI22D0BWP7T port map(A1 => gl_ram_n_240, A2 => gl_ram_n_44, B1 => gl_ram_n_242, B2 => gl_ram_n_32, ZN => gl_ram_n_293);
  gl_ram_g28597 : AOI22D0BWP7T port map(A1 => gl_ram_n_238, A2 => gl_ram_n_34, B1 => gl_ram_n_257, B2 => gl_ram_n_33, ZN => gl_ram_n_292);
  gl_ram_g28598 : AOI22D0BWP7T port map(A1 => gl_ram_n_255, A2 => gl_ram_n_44, B1 => gl_ram_n_243, B2 => gl_ram_n_32, ZN => gl_ram_n_291);
  gl_ram_g28599 : AOI22D0BWP7T port map(A1 => gl_ram_n_235, A2 => gl_ram_n_33, B1 => gl_ram_n_252, B2 => gl_ram_n_36, ZN => gl_ram_n_290);
  gl_ram_g28600 : AOI22D0BWP7T port map(A1 => gl_ram_n_237, A2 => gl_ram_n_34, B1 => gl_ram_n_239, B2 => gl_ram_n_33, ZN => gl_ram_n_289);
  gl_ram_g28601 : NR2XD0BWP7T port map(A1 => gl_ram_n_209, A2 => sig_logic_x(3), ZN => gl_ram_n_288);
  gl_ram_g28602 : FA1D0BWP7T port map(A => gl_ram_y_grid(1), B => gl_ram_x_grid(2), CI => gl_ram_n_16, CO => gl_ram_n_270, S => gl_ram_n_271);
  gl_ram_g28603 : ND4D0BWP7T port map(A1 => gl_ram_n_130, A2 => gl_ram_n_142, A3 => gl_ram_n_152, A4 => gl_ram_n_147, ZN => gl_ram_n_269);
  gl_ram_g28604 : ND4D0BWP7T port map(A1 => gl_ram_n_196, A2 => gl_ram_n_195, A3 => gl_ram_n_194, A4 => gl_ram_n_193, ZN => gl_ram_n_268);
  gl_ram_g28605 : ND4D0BWP7T port map(A1 => gl_ram_n_79, A2 => gl_ram_n_139, A3 => gl_ram_n_76, A4 => gl_ram_n_77, ZN => gl_ram_n_267);
  gl_ram_g28606 : ND4D0BWP7T port map(A1 => gl_ram_n_104, A2 => gl_ram_n_173, A3 => gl_ram_n_161, A4 => gl_ram_n_192, ZN => gl_ram_n_266);
  gl_ram_g28607 : ND4D0BWP7T port map(A1 => gl_ram_n_170, A2 => gl_ram_n_200, A3 => gl_ram_n_108, A4 => gl_ram_n_132, ZN => gl_ram_n_265);
  gl_ram_g28608 : ND4D0BWP7T port map(A1 => gl_ram_n_125, A2 => gl_ram_n_174, A3 => gl_ram_n_141, A4 => gl_ram_n_172, ZN => gl_ram_n_264);
  gl_ram_g28609 : ND4D0BWP7T port map(A1 => gl_ram_n_176, A2 => gl_ram_n_178, A3 => gl_ram_n_73, A4 => gl_ram_n_75, ZN => gl_ram_n_263);
  gl_ram_g28610 : ND4D0BWP7T port map(A1 => gl_ram_n_189, A2 => gl_ram_n_117, A3 => gl_ram_n_188, A4 => gl_ram_n_186, ZN => gl_ram_n_262);
  gl_ram_g28611 : ND4D0BWP7T port map(A1 => gl_ram_n_182, A2 => gl_ram_n_185, A3 => gl_ram_n_183, A4 => gl_ram_n_202, ZN => gl_ram_n_261);
  gl_ram_g28612 : ND4D0BWP7T port map(A1 => gl_ram_n_175, A2 => gl_ram_n_63, A3 => gl_ram_n_184, A4 => gl_ram_n_153, ZN => gl_ram_n_260);
  gl_ram_g28613 : NR2XD0BWP7T port map(A1 => gl_ram_n_231, A2 => gl_ram_n_207, ZN => gl_ram_n_287);
  gl_ram_g28614 : NR2XD0BWP7T port map(A1 => gl_ram_n_230, A2 => gl_ram_n_207, ZN => gl_ram_n_286);
  gl_ram_g28615 : NR2XD0BWP7T port map(A1 => gl_ram_n_231, A2 => gl_ram_n_205, ZN => gl_ram_n_285);
  gl_ram_g28616 : NR2XD0BWP7T port map(A1 => gl_ram_n_230, A2 => gl_ram_n_205, ZN => gl_ram_n_284);
  gl_ram_g28617 : NR2XD0BWP7T port map(A1 => gl_ram_n_231, A2 => gl_ram_n_208, ZN => gl_ram_n_283);
  gl_ram_g28618 : NR2XD0BWP7T port map(A1 => gl_ram_n_230, A2 => gl_ram_n_208, ZN => gl_ram_n_282);
  gl_ram_g28619 : NR2XD0BWP7T port map(A1 => gl_ram_n_231, A2 => gl_ram_n_206, ZN => gl_ram_n_281);
  gl_ram_g28620 : NR2XD0BWP7T port map(A1 => gl_ram_n_230, A2 => gl_ram_n_206, ZN => gl_ram_n_280);
  gl_ram_g28621 : NR2XD0BWP7T port map(A1 => gl_ram_n_232, A2 => gl_ram_n_207, ZN => gl_ram_n_279);
  gl_ram_g28622 : NR2XD0BWP7T port map(A1 => gl_ram_n_233, A2 => gl_ram_n_207, ZN => gl_ram_n_278);
  gl_ram_g28623 : NR2XD0BWP7T port map(A1 => gl_ram_n_233, A2 => gl_ram_n_206, ZN => gl_ram_n_277);
  gl_ram_g28624 : NR2XD0BWP7T port map(A1 => gl_ram_n_232, A2 => gl_ram_n_208, ZN => gl_ram_n_276);
  gl_ram_g28625 : NR2XD0BWP7T port map(A1 => gl_ram_n_232, A2 => gl_ram_n_206, ZN => gl_ram_n_275);
  gl_ram_g28626 : NR2XD0BWP7T port map(A1 => gl_ram_n_233, A2 => gl_ram_n_208, ZN => gl_ram_n_274);
  gl_ram_g28627 : NR2XD0BWP7T port map(A1 => gl_ram_n_232, A2 => gl_ram_n_205, ZN => gl_ram_n_273);
  gl_ram_g28628 : NR2XD0BWP7T port map(A1 => gl_ram_n_233, A2 => gl_ram_n_205, ZN => gl_ram_n_272);
  gl_ram_g28629 : ND4D0BWP7T port map(A1 => gl_ram_n_109, A2 => gl_ram_n_112, A3 => gl_ram_n_106, A4 => gl_ram_n_110, ZN => gl_ram_n_259);
  gl_ram_g28630 : ND4D0BWP7T port map(A1 => gl_ram_n_164, A2 => gl_ram_n_105, A3 => gl_ram_n_107, A4 => gl_ram_n_82, ZN => gl_ram_n_258);
  gl_ram_g28631 : ND4D0BWP7T port map(A1 => gl_ram_n_87, A2 => gl_ram_n_88, A3 => gl_ram_n_84, A4 => gl_ram_n_85, ZN => gl_ram_n_257);
  gl_ram_g28632 : ND4D0BWP7T port map(A1 => gl_ram_n_156, A2 => gl_ram_n_148, A3 => gl_ram_n_155, A4 => gl_ram_n_163, ZN => gl_ram_n_256);
  gl_ram_g28633 : ND4D0BWP7T port map(A1 => gl_ram_n_145, A2 => gl_ram_n_154, A3 => gl_ram_n_140, A4 => gl_ram_n_169, ZN => gl_ram_n_255);
  gl_ram_g28634 : ND4D0BWP7T port map(A1 => gl_ram_n_201, A2 => gl_ram_n_159, A3 => gl_ram_n_138, A4 => gl_ram_n_136, ZN => gl_ram_n_254);
  gl_ram_g28635 : ND4D0BWP7T port map(A1 => gl_ram_n_61, A2 => gl_ram_n_171, A3 => gl_ram_n_146, A4 => gl_ram_n_149, ZN => gl_ram_n_253);
  gl_ram_g28636 : ND4D0BWP7T port map(A1 => gl_ram_n_65, A2 => gl_ram_n_69, A3 => gl_ram_n_68, A4 => gl_ram_n_64, ZN => gl_ram_n_252);
  gl_ram_g28637 : ND4D0BWP7T port map(A1 => gl_ram_n_160, A2 => gl_ram_n_134, A3 => gl_ram_n_133, A4 => gl_ram_n_131, ZN => gl_ram_n_251);
  gl_ram_g28638 : ND4D0BWP7T port map(A1 => gl_ram_n_127, A2 => gl_ram_n_128, A3 => gl_ram_n_166, A4 => gl_ram_n_167, ZN => gl_ram_n_250);
  gl_ram_g28639 : ND4D0BWP7T port map(A1 => gl_ram_n_121, A2 => gl_ram_n_124, A3 => gl_ram_n_122, A4 => gl_ram_n_123, ZN => gl_ram_n_249);
  gl_ram_g28640 : ND4D0BWP7T port map(A1 => gl_ram_n_119, A2 => gl_ram_n_197, A3 => gl_ram_n_118, A4 => gl_ram_n_158, ZN => gl_ram_n_248);
  gl_ram_g28641 : ND4D0BWP7T port map(A1 => gl_ram_n_113, A2 => gl_ram_n_116, A3 => gl_ram_n_115, A4 => gl_ram_n_180, ZN => gl_ram_n_247);
  gl_ram_g28642 : ND4D0BWP7T port map(A1 => gl_ram_n_181, A2 => gl_ram_n_204, A3 => gl_ram_n_168, A4 => gl_ram_n_150, ZN => gl_ram_n_246);
  gl_ram_g28643 : ND4D0BWP7T port map(A1 => gl_ram_n_101, A2 => gl_ram_n_103, A3 => gl_ram_n_179, A4 => gl_ram_n_151, ZN => gl_ram_n_245);
  gl_ram_g28644 : ND4D0BWP7T port map(A1 => gl_ram_n_97, A2 => gl_ram_n_100, A3 => gl_ram_n_98, A4 => gl_ram_n_99, ZN => gl_ram_n_244);
  gl_ram_g28645 : ND4D0BWP7T port map(A1 => gl_ram_n_111, A2 => gl_ram_n_129, A3 => gl_ram_n_143, A4 => gl_ram_n_144, ZN => gl_ram_n_243);
  gl_ram_g28646 : ND4D0BWP7T port map(A1 => gl_ram_n_93, A2 => gl_ram_n_96, A3 => gl_ram_n_94, A4 => gl_ram_n_95, ZN => gl_ram_n_242);
  gl_ram_g28647 : ND4D0BWP7T port map(A1 => gl_ram_n_191, A2 => gl_ram_n_102, A3 => gl_ram_n_78, A4 => gl_ram_n_177, ZN => gl_ram_n_241);
  gl_ram_g28648 : ND4D0BWP7T port map(A1 => gl_ram_n_90, A2 => gl_ram_n_92, A3 => gl_ram_n_89, A4 => gl_ram_n_91, ZN => gl_ram_n_240);
  gl_ram_g28649 : ND4D0BWP7T port map(A1 => gl_ram_n_72, A2 => gl_ram_n_165, A3 => gl_ram_n_120, A4 => gl_ram_n_81, ZN => gl_ram_n_239);
  gl_ram_g28650 : ND4D0BWP7T port map(A1 => gl_ram_n_83, A2 => gl_ram_n_162, A3 => gl_ram_n_80, A4 => gl_ram_n_203, ZN => gl_ram_n_238);
  gl_ram_g28651 : ND4D0BWP7T port map(A1 => gl_ram_n_66, A2 => gl_ram_n_70, A3 => gl_ram_n_67, A4 => gl_ram_n_135, ZN => gl_ram_n_237);
  gl_ram_g28652 : ND4D0BWP7T port map(A1 => gl_ram_n_74, A2 => gl_ram_n_114, A3 => gl_ram_n_126, A4 => gl_ram_n_71, ZN => gl_ram_n_236);
  gl_ram_g28653 : ND4D0BWP7T port map(A1 => gl_ram_n_157, A2 => gl_ram_n_137, A3 => gl_ram_n_62, A4 => gl_ram_n_198, ZN => gl_ram_n_235);
  gl_ram_g28654 : ND4D0BWP7T port map(A1 => gl_ram_n_86, A2 => gl_ram_n_199, A3 => gl_ram_n_187, A4 => gl_ram_n_190, ZN => gl_ram_n_234);
  gl_ram_g28655 : NR2D1BWP7T port map(A1 => gl_ram_n_213, A2 => sig_middelsteknop, ZN => gl_ram_n_233);
  gl_ram_g28656 : AN2D1BWP7T port map(A1 => gl_ram_n_212, A2 => gl_ram_n_6, Z => gl_ram_n_232);
  gl_ram_g28657 : NR2XD0BWP7T port map(A1 => gl_ram_n_214, A2 => sig_middelsteknop, ZN => gl_ram_n_231);
  gl_ram_g28658 : NR2XD0BWP7T port map(A1 => gl_ram_n_211, A2 => sig_middelsteknop, ZN => gl_ram_n_230);
  gl_ram_g28659 : CKAN2D1BWP7T port map(A1 => gl_ram_n_214, A2 => gl_ram_n_46, Z => gl_ram_n_229);
  gl_ram_g28660 : NR2XD0BWP7T port map(A1 => gl_ram_n_210, A2 => gl_ram_n_42, ZN => gl_ram_n_228);
  gl_ram_g28661 : CKAN2D1BWP7T port map(A1 => gl_ram_n_214, A2 => gl_ram_n_43, Z => gl_ram_n_227);
  gl_ram_g28662 : NR2XD0BWP7T port map(A1 => gl_ram_n_212, A2 => gl_ram_n_47, ZN => gl_ram_n_226);
  gl_ram_g28663 : NR2XD0BWP7T port map(A1 => gl_ram_n_212, A2 => gl_ram_n_42, ZN => gl_ram_n_225);
  gl_ram_g28664 : AOI22D0BWP7T port map(A1 => gl_ram_n_58, A2 => gl_ram_ram_96(2), B1 => gl_ram_n_53, B2 => gl_ram_ram_99(2), ZN => gl_ram_n_221);
  gl_ram_g28665 : OA21D0BWP7T port map(A1 => gl_ram_n_19, A2 => gl_ram_n_5, B => gl_ram_n_209, Z => gl_ram_n_220);
  gl_ram_g28666 : AOI22D0BWP7T port map(A1 => gl_ram_n_58, A2 => gl_ram_ram_96(1), B1 => gl_ram_n_53, B2 => gl_ram_ram_99(1), ZN => gl_ram_n_219);
  gl_ram_g28667 : AOI22D0BWP7T port map(A1 => gl_ram_n_52, A2 => gl_ram_ram_97(1), B1 => gl_ram_n_51, B2 => gl_ram_ram_98(1), ZN => gl_ram_n_218);
  gl_ram_g28668 : AOI22D0BWP7T port map(A1 => gl_ram_n_58, A2 => gl_ram_ram_96(0), B1 => gl_ram_n_53, B2 => gl_ram_ram_99(0), ZN => gl_ram_n_217);
  gl_ram_g28669 : AOI22D0BWP7T port map(A1 => gl_ram_n_52, A2 => gl_ram_ram_97(2), B1 => gl_ram_n_51, B2 => gl_ram_ram_98(2), ZN => gl_ram_n_216);
  gl_ram_g28670 : AOI22D0BWP7T port map(A1 => gl_ram_n_52, A2 => gl_ram_ram_97(0), B1 => gl_ram_n_51, B2 => gl_ram_ram_98(0), ZN => gl_ram_n_215);
  gl_ram_g28671 : NR2XD0BWP7T port map(A1 => gl_ram_n_210, A2 => gl_ram_n_47, ZN => gl_ram_n_224);
  gl_ram_g28672 : CKAN2D1BWP7T port map(A1 => gl_ram_n_213, A2 => gl_ram_n_43, Z => gl_ram_n_223);
  gl_ram_g28673 : CKAN2D1BWP7T port map(A1 => gl_ram_n_213, A2 => gl_ram_n_46, Z => gl_ram_n_222);
  gl_ram_g28674 : INVD0BWP7T port map(I => gl_ram_n_210, ZN => gl_ram_n_211);
  gl_ram_g28675 : AOI22D0BWP7T port map(A1 => gl_ram_n_40, A2 => gl_ram_ram_21(2), B1 => gl_ram_n_39, B2 => gl_ram_ram_19(2), ZN => gl_ram_n_204);
  gl_ram_g28676 : AOI22D0BWP7T port map(A1 => gl_ram_n_38, A2 => gl_ram_ram_72(2), B1 => gl_ram_n_29, B2 => gl_ram_ram_79(2), ZN => gl_ram_n_203);
  gl_ram_g28677 : AOI22D0BWP7T port map(A1 => gl_ram_n_30, A2 => gl_ram_ram_65(0), B1 => gl_ram_n_29, B2 => gl_ram_ram_71(0), ZN => gl_ram_n_202);
  gl_ram_g28678 : AOI22D0BWP7T port map(A1 => gl_ram_n_28, A2 => gl_ram_ram_90(1), B1 => gl_ram_n_31, B2 => gl_ram_ram_94(1), ZN => gl_ram_n_201);
  gl_ram_g28679 : AOI22D0BWP7T port map(A1 => gl_ram_n_40, A2 => gl_ram_ram_53(0), B1 => gl_ram_n_39, B2 => gl_ram_ram_51(0), ZN => gl_ram_n_200);
  gl_ram_g28680 : AOI22D0BWP7T port map(A1 => gl_ram_n_40, A2 => gl_ram_ram_85(0), B1 => gl_ram_n_39, B2 => gl_ram_ram_83(0), ZN => gl_ram_n_199);
  gl_ram_g28681 : AOI22D0BWP7T port map(A1 => gl_ram_n_38, A2 => gl_ram_ram_24(2), B1 => gl_ram_n_31, B2 => gl_ram_ram_30(2), ZN => gl_ram_n_198);
  gl_ram_g28682 : AOI22D0BWP7T port map(A1 => gl_ram_n_40, A2 => gl_ram_ram_29(1), B1 => gl_ram_n_39, B2 => gl_ram_ram_27(1), ZN => gl_ram_n_197);
  gl_ram_g28683 : AOI22D0BWP7T port map(A1 => gl_ram_n_28, A2 => gl_ram_ram_50(2), B1 => gl_ram_n_31, B2 => gl_ram_ram_54(2), ZN => gl_ram_n_196);
  gl_ram_g28684 : AOI22D0BWP7T port map(A1 => gl_ram_n_40, A2 => gl_ram_ram_53(2), B1 => gl_ram_n_39, B2 => gl_ram_ram_51(2), ZN => gl_ram_n_195);
  gl_ram_g28685 : AOI22D0BWP7T port map(A1 => gl_ram_n_30, A2 => gl_ram_ram_49(2), B1 => gl_ram_n_29, B2 => gl_ram_ram_55(2), ZN => gl_ram_n_194);
  gl_ram_g28686 : AOI22D0BWP7T port map(A1 => gl_ram_n_38, A2 => gl_ram_ram_48(2), B1 => gl_ram_n_41, B2 => gl_ram_ram_52(2), ZN => gl_ram_n_193);
  gl_ram_g28687 : AOI22D0BWP7T port map(A1 => gl_ram_n_38, A2 => gl_ram_ram_56(0), B1 => gl_ram_n_41, B2 => gl_ram_ram_60(0), ZN => gl_ram_n_192);
  gl_ram_g28688 : AOI22D0BWP7T port map(A1 => gl_ram_n_28, A2 => gl_ram_ram_34(2), B1 => gl_ram_n_31, B2 => gl_ram_ram_38(2), ZN => gl_ram_n_191);
  gl_ram_g28689 : AOI22D0BWP7T port map(A1 => gl_ram_n_30, A2 => gl_ram_ram_81(0), B1 => gl_ram_n_29, B2 => gl_ram_ram_87(0), ZN => gl_ram_n_190);
  gl_ram_g28690 : AOI22D0BWP7T port map(A1 => gl_ram_n_40, A2 => gl_ram_ram_45(2), B1 => gl_ram_n_39, B2 => gl_ram_ram_43(2), ZN => gl_ram_n_189);
  gl_ram_g28691 : AOI22D0BWP7T port map(A1 => gl_ram_n_30, A2 => gl_ram_ram_41(2), B1 => gl_ram_n_29, B2 => gl_ram_ram_47(2), ZN => gl_ram_n_188);
  gl_ram_g28692 : AOI22D0BWP7T port map(A1 => gl_ram_n_41, A2 => gl_ram_ram_84(0), B1 => gl_ram_n_28, B2 => gl_ram_ram_82(0), ZN => gl_ram_n_187);
  gl_ram_g28693 : AOI22D0BWP7T port map(A1 => gl_ram_n_38, A2 => gl_ram_ram_40(2), B1 => gl_ram_n_31, B2 => gl_ram_ram_46(2), ZN => gl_ram_n_186);
  gl_ram_g28694 : AOI22D0BWP7T port map(A1 => gl_ram_n_40, A2 => gl_ram_ram_69(0), B1 => gl_ram_n_39, B2 => gl_ram_ram_67(0), ZN => gl_ram_n_185);
  gl_ram_g28695 : AOI22D0BWP7T port map(A1 => gl_ram_n_30, A2 => gl_ram_ram_9(2), B1 => gl_ram_n_29, B2 => gl_ram_ram_15(2), ZN => gl_ram_n_184);
  gl_ram_g28696 : AOI22D0BWP7T port map(A1 => gl_ram_n_41, A2 => gl_ram_ram_68(0), B1 => gl_ram_n_28, B2 => gl_ram_ram_66(0), ZN => gl_ram_n_183);
  gl_ram_g28697 : AOI22D0BWP7T port map(A1 => gl_ram_n_38, A2 => gl_ram_ram_64(0), B1 => gl_ram_n_31, B2 => gl_ram_ram_70(0), ZN => gl_ram_n_182);
  gl_ram_g28698 : AOI22D0BWP7T port map(A1 => gl_ram_n_28, A2 => gl_ram_ram_18(2), B1 => gl_ram_n_31, B2 => gl_ram_ram_22(2), ZN => gl_ram_n_181);
  gl_ram_g28699 : AOI22D0BWP7T port map(A1 => gl_ram_n_30, A2 => gl_ram_ram_9(1), B1 => gl_ram_n_29, B2 => gl_ram_ram_15(1), ZN => gl_ram_n_180);
  gl_ram_g28700 : AOI22D0BWP7T port map(A1 => gl_ram_n_41, A2 => gl_ram_ram_44(1), B1 => gl_ram_n_28, B2 => gl_ram_ram_42(1), ZN => gl_ram_n_179);
  gl_ram_g28701 : AOI22D0BWP7T port map(A1 => gl_ram_n_40, A2 => gl_ram_ram_45(0), B1 => gl_ram_n_39, B2 => gl_ram_ram_43(0), ZN => gl_ram_n_178);
  gl_ram_g28702 : AOI22D0BWP7T port map(A1 => gl_ram_n_38, A2 => gl_ram_ram_32(2), B1 => gl_ram_n_41, B2 => gl_ram_ram_36(2), ZN => gl_ram_n_177);
  gl_ram_g28703 : AOI22D0BWP7T port map(A1 => gl_ram_n_28, A2 => gl_ram_ram_42(0), B1 => gl_ram_n_31, B2 => gl_ram_ram_46(0), ZN => gl_ram_n_176);
  gl_ram_g28704 : AOI22D0BWP7T port map(A1 => gl_ram_n_28, A2 => gl_ram_ram_10(2), B1 => gl_ram_n_31, B2 => gl_ram_ram_14(2), ZN => gl_ram_n_175);
  gl_ram_g28705 : AOI22D0BWP7T port map(A1 => gl_ram_n_41, A2 => gl_ram_ram_4(2), B1 => gl_ram_n_28, B2 => gl_ram_ram_2(2), ZN => gl_ram_n_174);
  gl_ram_g28706 : AOI22D0BWP7T port map(A1 => gl_ram_n_40, A2 => gl_ram_ram_61(0), B1 => gl_ram_n_39, B2 => gl_ram_ram_59(0), ZN => gl_ram_n_173);
  gl_ram_g28707 : AOI22D0BWP7T port map(A1 => gl_ram_n_38, A2 => gl_ram_ram_0(2), B1 => gl_ram_n_31, B2 => gl_ram_ram_6(2), ZN => gl_ram_n_172);
  gl_ram_g28708 : AOI22D0BWP7T port map(A1 => gl_ram_n_40, A2 => gl_ram_ram_77(1), B1 => gl_ram_n_39, B2 => gl_ram_ram_75(1), ZN => gl_ram_n_171);
  gl_ram_g28709 : AOI22D0BWP7T port map(A1 => gl_ram_n_28, A2 => gl_ram_ram_50(0), B1 => gl_ram_n_31, B2 => gl_ram_ram_54(0), ZN => gl_ram_n_170);
  gl_ram_g28710 : AOI22D0BWP7T port map(A1 => gl_ram_n_38, A2 => gl_ram_ram_0(0), B1 => gl_ram_n_31, B2 => gl_ram_ram_6(0), ZN => gl_ram_n_169);
  gl_ram_g28711 : AOI22D0BWP7T port map(A1 => gl_ram_n_30, A2 => gl_ram_ram_17(2), B1 => gl_ram_n_29, B2 => gl_ram_ram_23(2), ZN => gl_ram_n_168);
  gl_ram_g28712 : AOI22D0BWP7T port map(A1 => gl_ram_n_38, A2 => gl_ram_ram_64(1), B1 => gl_ram_n_41, B2 => gl_ram_ram_68(1), ZN => gl_ram_n_167);
  gl_ram_g28713 : AOI22D0BWP7T port map(A1 => gl_ram_n_30, A2 => gl_ram_ram_65(1), B1 => gl_ram_n_29, B2 => gl_ram_ram_71(1), ZN => gl_ram_n_166);
  gl_ram_g28714 : AOI22D0BWP7T port map(A1 => gl_ram_n_40, A2 => gl_ram_ram_93(0), B1 => gl_ram_n_39, B2 => gl_ram_ram_91(0), ZN => gl_ram_n_165);
  gl_ram_g28715 : AOI22D0BWP7T port map(A1 => gl_ram_n_28, A2 => gl_ram_ram_26(0), B1 => gl_ram_n_31, B2 => gl_ram_ram_30(0), ZN => gl_ram_n_164);
  gl_ram_g28716 : AOI22D0BWP7T port map(A1 => gl_ram_n_38, A2 => gl_ram_ram_16(0), B1 => gl_ram_n_31, B2 => gl_ram_ram_22(0), ZN => gl_ram_n_163);
  gl_ram_g28717 : AOI22D0BWP7T port map(A1 => gl_ram_n_40, A2 => gl_ram_ram_77(2), B1 => gl_ram_n_39, B2 => gl_ram_ram_75(2), ZN => gl_ram_n_162);
  gl_ram_g28718 : AOI22D0BWP7T port map(A1 => gl_ram_n_30, A2 => gl_ram_ram_57(0), B1 => gl_ram_n_29, B2 => gl_ram_ram_63(0), ZN => gl_ram_n_161);
  gl_ram_g28719 : AOI22D0BWP7T port map(A1 => gl_ram_n_28, A2 => gl_ram_ram_82(1), B1 => gl_ram_n_31, B2 => gl_ram_ram_86(1), ZN => gl_ram_n_160);
  gl_ram_g28720 : AOI22D0BWP7T port map(A1 => gl_ram_n_40, A2 => gl_ram_ram_93(1), B1 => gl_ram_n_39, B2 => gl_ram_ram_91(1), ZN => gl_ram_n_159);
  gl_ram_g28721 : AOI22D0BWP7T port map(A1 => gl_ram_n_30, A2 => gl_ram_ram_25(1), B1 => gl_ram_n_29, B2 => gl_ram_ram_31(1), ZN => gl_ram_n_158);
  gl_ram_g28722 : AOI22D0BWP7T port map(A1 => gl_ram_n_40, A2 => gl_ram_ram_29(2), B1 => gl_ram_n_39, B2 => gl_ram_ram_27(2), ZN => gl_ram_n_157);
  gl_ram_g28723 : AOI22D0BWP7T port map(A1 => gl_ram_n_40, A2 => gl_ram_ram_21(0), B1 => gl_ram_n_39, B2 => gl_ram_ram_19(0), ZN => gl_ram_n_156);
  gl_ram_g28724 : AOI22D0BWP7T port map(A1 => gl_ram_n_30, A2 => gl_ram_ram_17(0), B1 => gl_ram_n_29, B2 => gl_ram_ram_23(0), ZN => gl_ram_n_155);
  gl_ram_g28725 : AOI22D0BWP7T port map(A1 => gl_ram_n_41, A2 => gl_ram_ram_4(0), B1 => gl_ram_n_28, B2 => gl_ram_ram_2(0), ZN => gl_ram_n_154);
  gl_ram_g28726 : AOI22D0BWP7T port map(A1 => gl_ram_n_38, A2 => gl_ram_ram_8(2), B1 => gl_ram_n_41, B2 => gl_ram_ram_12(2), ZN => gl_ram_n_153);
  gl_ram_g28727 : AOI22D0BWP7T port map(A1 => gl_ram_n_30, A2 => gl_ram_ram_9(0), B1 => gl_ram_n_29, B2 => gl_ram_ram_15(0), ZN => gl_ram_n_152);
  gl_ram_g28728 : AOI22D0BWP7T port map(A1 => gl_ram_n_30, A2 => gl_ram_ram_41(1), B1 => gl_ram_n_29, B2 => gl_ram_ram_47(1), ZN => gl_ram_n_151);
  gl_ram_g28729 : AOI22D0BWP7T port map(A1 => gl_ram_n_38, A2 => gl_ram_ram_16(2), B1 => gl_ram_n_41, B2 => gl_ram_ram_20(2), ZN => gl_ram_n_150);
  gl_ram_g28730 : AOI22D0BWP7T port map(A1 => gl_ram_n_38, A2 => gl_ram_ram_72(1), B1 => gl_ram_n_41, B2 => gl_ram_ram_76(1), ZN => gl_ram_n_149);
  gl_ram_g28731 : AOI22D0BWP7T port map(A1 => gl_ram_n_41, A2 => gl_ram_ram_20(0), B1 => gl_ram_n_28, B2 => gl_ram_ram_18(0), ZN => gl_ram_n_148);
  gl_ram_g28732 : AOI22D0BWP7T port map(A1 => gl_ram_n_38, A2 => gl_ram_ram_8(0), B1 => gl_ram_n_31, B2 => gl_ram_ram_14(0), ZN => gl_ram_n_147);
  gl_ram_g28733 : AOI22D0BWP7T port map(A1 => gl_ram_n_30, A2 => gl_ram_ram_73(1), B1 => gl_ram_n_29, B2 => gl_ram_ram_79(1), ZN => gl_ram_n_146);
  gl_ram_g28734 : AOI22D0BWP7T port map(A1 => gl_ram_n_40, A2 => gl_ram_ram_5(0), B1 => gl_ram_n_39, B2 => gl_ram_ram_3(0), ZN => gl_ram_n_145);
  gl_ram_g28735 : AOI22D0BWP7T port map(A1 => gl_ram_n_38, A2 => gl_ram_ram_32(0), B1 => gl_ram_n_31, B2 => gl_ram_ram_38(0), ZN => gl_ram_n_144);
  gl_ram_g28736 : AOI22D0BWP7T port map(A1 => gl_ram_n_30, A2 => gl_ram_ram_33(0), B1 => gl_ram_n_29, B2 => gl_ram_ram_39(0), ZN => gl_ram_n_143);
  gl_ram_g28737 : AOI22D0BWP7T port map(A1 => gl_ram_n_41, A2 => gl_ram_ram_12(0), B1 => gl_ram_n_28, B2 => gl_ram_ram_10(0), ZN => gl_ram_n_142);
  gl_ram_g28738 : AOI22D0BWP7T port map(A1 => gl_ram_n_30, A2 => gl_ram_ram_1(2), B1 => gl_ram_n_29, B2 => gl_ram_ram_7(2), ZN => gl_ram_n_141);
  gl_ram_g28739 : AOI22D0BWP7T port map(A1 => gl_ram_n_30, A2 => gl_ram_ram_1(0), B1 => gl_ram_n_29, B2 => gl_ram_ram_7(0), ZN => gl_ram_n_140);
  gl_ram_g28740 : AOI22D0BWP7T port map(A1 => gl_ram_n_40, A2 => gl_ram_ram_85(2), B1 => gl_ram_n_39, B2 => gl_ram_ram_83(2), ZN => gl_ram_n_139);
  gl_ram_g28741 : AOI22D0BWP7T port map(A1 => gl_ram_n_30, A2 => gl_ram_ram_89(1), B1 => gl_ram_n_29, B2 => gl_ram_ram_95(1), ZN => gl_ram_n_138);
  gl_ram_g28742 : NR2XD0BWP7T port map(A1 => gl_ram_n_60, A2 => gl_ram_ram_position(1), ZN => gl_ram_n_214);
  gl_ram_g28743 : INR2XD0BWP7T port map(A1 => gl_ram_n_59, B1 => gl_ram_ram_position(1), ZN => gl_ram_n_213);
  gl_ram_g28744 : ND2D1BWP7T port map(A1 => gl_ram_n_59, A2 => gl_ram_ram_position(1), ZN => gl_ram_n_212);
  gl_ram_g28745 : IND2D1BWP7T port map(A1 => gl_ram_n_60, B1 => gl_ram_ram_position(1), ZN => gl_ram_n_210);
  gl_ram_g28746 : ND2D1BWP7T port map(A1 => gl_ram_n_19, A2 => gl_ram_n_5, ZN => gl_ram_n_209);
  gl_ram_g28747 : AOI21D0BWP7T port map(A1 => gl_ram_n_43, A2 => gl_ram_ram_position(0), B => sig_middelsteknop, ZN => gl_ram_n_208);
  gl_ram_g28748 : AOI21D0BWP7T port map(A1 => gl_ram_n_46, A2 => gl_ram_n_3, B => sig_middelsteknop, ZN => gl_ram_n_207);
  gl_ram_g28749 : AOI21D0BWP7T port map(A1 => gl_ram_n_43, A2 => gl_ram_n_3, B => sig_middelsteknop, ZN => gl_ram_n_206);
  gl_ram_g28750 : AOI21D0BWP7T port map(A1 => gl_ram_n_46, A2 => gl_ram_ram_position(0), B => sig_middelsteknop, ZN => gl_ram_n_205);
  gl_ram_g28751 : AOI22D0BWP7T port map(A1 => gl_ram_n_41, A2 => gl_ram_ram_28(2), B1 => gl_ram_n_28, B2 => gl_ram_ram_26(2), ZN => gl_ram_n_137);
  gl_ram_g28752 : AOI22D0BWP7T port map(A1 => gl_ram_n_38, A2 => gl_ram_ram_88(1), B1 => gl_ram_n_41, B2 => gl_ram_ram_92(1), ZN => gl_ram_n_136);
  gl_ram_g28753 : AOI22D0BWP7T port map(A1 => gl_ram_n_30, A2 => gl_ram_ram_73(0), B1 => gl_ram_n_29, B2 => gl_ram_ram_79(0), ZN => gl_ram_n_135);
  gl_ram_g28754 : AOI22D0BWP7T port map(A1 => gl_ram_n_40, A2 => gl_ram_ram_85(1), B1 => gl_ram_n_39, B2 => gl_ram_ram_83(1), ZN => gl_ram_n_134);
  gl_ram_g28755 : AOI22D0BWP7T port map(A1 => gl_ram_n_30, A2 => gl_ram_ram_81(1), B1 => gl_ram_n_29, B2 => gl_ram_ram_87(1), ZN => gl_ram_n_133);
  gl_ram_g28756 : AOI22D0BWP7T port map(A1 => gl_ram_n_38, A2 => gl_ram_ram_48(0), B1 => gl_ram_n_29, B2 => gl_ram_ram_55(0), ZN => gl_ram_n_132);
  gl_ram_g28757 : AOI22D0BWP7T port map(A1 => gl_ram_n_38, A2 => gl_ram_ram_80(1), B1 => gl_ram_n_41, B2 => gl_ram_ram_84(1), ZN => gl_ram_n_131);
  gl_ram_g28758 : AOI22D0BWP7T port map(A1 => gl_ram_n_40, A2 => gl_ram_ram_13(0), B1 => gl_ram_n_39, B2 => gl_ram_ram_11(0), ZN => gl_ram_n_130);
  gl_ram_g28759 : AOI22D0BWP7T port map(A1 => gl_ram_n_41, A2 => gl_ram_ram_36(0), B1 => gl_ram_n_28, B2 => gl_ram_ram_34(0), ZN => gl_ram_n_129);
  gl_ram_g28760 : AOI22D0BWP7T port map(A1 => gl_ram_n_40, A2 => gl_ram_ram_69(1), B1 => gl_ram_n_39, B2 => gl_ram_ram_67(1), ZN => gl_ram_n_128);
  gl_ram_g28761 : AOI22D0BWP7T port map(A1 => gl_ram_n_28, A2 => gl_ram_ram_66(1), B1 => gl_ram_n_31, B2 => gl_ram_ram_70(1), ZN => gl_ram_n_127);
  gl_ram_g28762 : AOI22D0BWP7T port map(A1 => gl_ram_n_41, A2 => gl_ram_ram_68(2), B1 => gl_ram_n_30, B2 => gl_ram_ram_65(2), ZN => gl_ram_n_126);
  gl_ram_g28763 : AOI22D0BWP7T port map(A1 => gl_ram_n_40, A2 => gl_ram_ram_5(2), B1 => gl_ram_n_39, B2 => gl_ram_ram_3(2), ZN => gl_ram_n_125);
  gl_ram_g28764 : AOI22D0BWP7T port map(A1 => gl_ram_n_40, A2 => gl_ram_ram_61(1), B1 => gl_ram_n_39, B2 => gl_ram_ram_59(1), ZN => gl_ram_n_124);
  gl_ram_g28765 : AOI22D0BWP7T port map(A1 => gl_ram_n_30, A2 => gl_ram_ram_57(1), B1 => gl_ram_n_29, B2 => gl_ram_ram_63(1), ZN => gl_ram_n_123);
  gl_ram_g28766 : AOI22D0BWP7T port map(A1 => gl_ram_n_41, A2 => gl_ram_ram_60(1), B1 => gl_ram_n_28, B2 => gl_ram_ram_58(1), ZN => gl_ram_n_122);
  gl_ram_g28767 : AOI22D0BWP7T port map(A1 => gl_ram_n_38, A2 => gl_ram_ram_56(1), B1 => gl_ram_n_31, B2 => gl_ram_ram_62(1), ZN => gl_ram_n_121);
  gl_ram_g28768 : AOI22D0BWP7T port map(A1 => gl_ram_n_38, A2 => gl_ram_ram_88(0), B1 => gl_ram_n_41, B2 => gl_ram_ram_92(0), ZN => gl_ram_n_120);
  gl_ram_g28769 : AOI22D0BWP7T port map(A1 => gl_ram_n_28, A2 => gl_ram_ram_26(1), B1 => gl_ram_n_31, B2 => gl_ram_ram_30(1), ZN => gl_ram_n_119);
  gl_ram_g28770 : AOI22D0BWP7T port map(A1 => gl_ram_n_38, A2 => gl_ram_ram_24(1), B1 => gl_ram_n_41, B2 => gl_ram_ram_28(1), ZN => gl_ram_n_118);
  gl_ram_g28771 : AOI22D0BWP7T port map(A1 => gl_ram_n_41, A2 => gl_ram_ram_44(2), B1 => gl_ram_n_28, B2 => gl_ram_ram_42(2), ZN => gl_ram_n_117);
  gl_ram_g28772 : AOI22D0BWP7T port map(A1 => gl_ram_n_40, A2 => gl_ram_ram_13(1), B1 => gl_ram_n_39, B2 => gl_ram_ram_11(1), ZN => gl_ram_n_116);
  gl_ram_g28773 : AOI22D0BWP7T port map(A1 => gl_ram_n_41, A2 => gl_ram_ram_12(1), B1 => gl_ram_n_28, B2 => gl_ram_ram_10(1), ZN => gl_ram_n_115);
  gl_ram_g28774 : AOI22D0BWP7T port map(A1 => gl_ram_n_40, A2 => gl_ram_ram_69(2), B1 => gl_ram_n_39, B2 => gl_ram_ram_67(2), ZN => gl_ram_n_114);
  gl_ram_g28775 : AOI22D0BWP7T port map(A1 => gl_ram_n_38, A2 => gl_ram_ram_8(1), B1 => gl_ram_n_31, B2 => gl_ram_ram_14(1), ZN => gl_ram_n_113);
  gl_ram_g28776 : AOI22D0BWP7T port map(A1 => gl_ram_n_40, A2 => gl_ram_ram_21(1), B1 => gl_ram_n_39, B2 => gl_ram_ram_19(1), ZN => gl_ram_n_112);
  gl_ram_g28777 : AOI22D0BWP7T port map(A1 => gl_ram_n_40, A2 => gl_ram_ram_37(0), B1 => gl_ram_n_39, B2 => gl_ram_ram_35(0), ZN => gl_ram_n_111);
  gl_ram_g28778 : AOI22D0BWP7T port map(A1 => gl_ram_n_30, A2 => gl_ram_ram_17(1), B1 => gl_ram_n_29, B2 => gl_ram_ram_23(1), ZN => gl_ram_n_110);
  gl_ram_g28779 : AOI22D0BWP7T port map(A1 => gl_ram_n_28, A2 => gl_ram_ram_18(1), B1 => gl_ram_n_31, B2 => gl_ram_ram_22(1), ZN => gl_ram_n_109);
  gl_ram_g28780 : AOI22D0BWP7T port map(A1 => gl_ram_n_41, A2 => gl_ram_ram_52(0), B1 => gl_ram_n_30, B2 => gl_ram_ram_49(0), ZN => gl_ram_n_108);
  gl_ram_g28781 : AOI22D0BWP7T port map(A1 => gl_ram_n_38, A2 => gl_ram_ram_24(0), B1 => gl_ram_n_40, B2 => gl_ram_ram_29(0), ZN => gl_ram_n_107);
  gl_ram_g28782 : AOI22D0BWP7T port map(A1 => gl_ram_n_38, A2 => gl_ram_ram_16(1), B1 => gl_ram_n_41, B2 => gl_ram_ram_20(1), ZN => gl_ram_n_106);
  gl_ram_g28783 : AOI22D0BWP7T port map(A1 => gl_ram_n_30, A2 => gl_ram_ram_25(0), B1 => gl_ram_n_29, B2 => gl_ram_ram_31(0), ZN => gl_ram_n_105);
  gl_ram_g28784 : AOI22D0BWP7T port map(A1 => gl_ram_n_28, A2 => gl_ram_ram_58(0), B1 => gl_ram_n_31, B2 => gl_ram_ram_62(0), ZN => gl_ram_n_104);
  gl_ram_g28785 : AOI22D0BWP7T port map(A1 => gl_ram_n_40, A2 => gl_ram_ram_45(1), B1 => gl_ram_n_39, B2 => gl_ram_ram_43(1), ZN => gl_ram_n_103);
  gl_ram_g28786 : AOI22D0BWP7T port map(A1 => gl_ram_n_40, A2 => gl_ram_ram_37(2), B1 => gl_ram_n_39, B2 => gl_ram_ram_35(2), ZN => gl_ram_n_102);
  gl_ram_g28787 : AOI22D0BWP7T port map(A1 => gl_ram_n_38, A2 => gl_ram_ram_40(1), B1 => gl_ram_n_31, B2 => gl_ram_ram_46(1), ZN => gl_ram_n_101);
  gl_ram_g28788 : AOI22D0BWP7T port map(A1 => gl_ram_n_40, A2 => gl_ram_ram_53(1), B1 => gl_ram_n_39, B2 => gl_ram_ram_51(1), ZN => gl_ram_n_100);
  gl_ram_g28789 : AOI22D0BWP7T port map(A1 => gl_ram_n_30, A2 => gl_ram_ram_49(1), B1 => gl_ram_n_29, B2 => gl_ram_ram_55(1), ZN => gl_ram_n_99);
  gl_ram_g28790 : AOI22D0BWP7T port map(A1 => gl_ram_n_41, A2 => gl_ram_ram_52(1), B1 => gl_ram_n_28, B2 => gl_ram_ram_50(1), ZN => gl_ram_n_98);
  gl_ram_g28791 : AOI22D0BWP7T port map(A1 => gl_ram_n_38, A2 => gl_ram_ram_48(1), B1 => gl_ram_n_31, B2 => gl_ram_ram_54(1), ZN => gl_ram_n_97);
  gl_ram_g28792 : AOI22D0BWP7T port map(A1 => gl_ram_n_40, A2 => gl_ram_ram_37(1), B1 => gl_ram_n_39, B2 => gl_ram_ram_35(1), ZN => gl_ram_n_96);
  gl_ram_g28793 : AOI22D0BWP7T port map(A1 => gl_ram_n_30, A2 => gl_ram_ram_33(1), B1 => gl_ram_n_29, B2 => gl_ram_ram_39(1), ZN => gl_ram_n_95);
  gl_ram_g28794 : AOI22D0BWP7T port map(A1 => gl_ram_n_41, A2 => gl_ram_ram_36(1), B1 => gl_ram_n_28, B2 => gl_ram_ram_34(1), ZN => gl_ram_n_94);
  gl_ram_g28795 : AOI22D0BWP7T port map(A1 => gl_ram_n_38, A2 => gl_ram_ram_32(1), B1 => gl_ram_n_31, B2 => gl_ram_ram_38(1), ZN => gl_ram_n_93);
  gl_ram_g28796 : AOI22D0BWP7T port map(A1 => gl_ram_n_40, A2 => gl_ram_ram_5(1), B1 => gl_ram_n_39, B2 => gl_ram_ram_3(1), ZN => gl_ram_n_92);
  gl_ram_g28797 : AOI22D0BWP7T port map(A1 => gl_ram_n_30, A2 => gl_ram_ram_1(1), B1 => gl_ram_n_29, B2 => gl_ram_ram_7(1), ZN => gl_ram_n_91);
  gl_ram_g28798 : AOI22D0BWP7T port map(A1 => gl_ram_n_28, A2 => gl_ram_ram_2(1), B1 => gl_ram_n_31, B2 => gl_ram_ram_6(1), ZN => gl_ram_n_90);
  gl_ram_g28799 : AOI22D0BWP7T port map(A1 => gl_ram_n_38, A2 => gl_ram_ram_0(1), B1 => gl_ram_n_41, B2 => gl_ram_ram_4(1), ZN => gl_ram_n_89);
  gl_ram_g28800 : AOI22D0BWP7T port map(A1 => gl_ram_n_30, A2 => gl_ram_ram_89(2), B1 => gl_ram_n_29, B2 => gl_ram_ram_95(2), ZN => gl_ram_n_88);
  gl_ram_g28801 : AOI22D0BWP7T port map(A1 => gl_ram_n_28, A2 => gl_ram_ram_90(2), B1 => gl_ram_n_31, B2 => gl_ram_ram_94(2), ZN => gl_ram_n_87);
  gl_ram_g28802 : AOI22D0BWP7T port map(A1 => gl_ram_n_38, A2 => gl_ram_ram_80(0), B1 => gl_ram_n_31, B2 => gl_ram_ram_86(0), ZN => gl_ram_n_86);
  gl_ram_g28803 : AOI22D0BWP7T port map(A1 => gl_ram_n_40, A2 => gl_ram_ram_93(2), B1 => gl_ram_n_39, B2 => gl_ram_ram_91(2), ZN => gl_ram_n_85);
  gl_ram_g28804 : AOI22D0BWP7T port map(A1 => gl_ram_n_38, A2 => gl_ram_ram_88(2), B1 => gl_ram_n_41, B2 => gl_ram_ram_92(2), ZN => gl_ram_n_84);
  gl_ram_g28805 : AOI22D0BWP7T port map(A1 => gl_ram_n_28, A2 => gl_ram_ram_74(2), B1 => gl_ram_n_31, B2 => gl_ram_ram_78(2), ZN => gl_ram_n_83);
  gl_ram_g28806 : AOI22D0BWP7T port map(A1 => gl_ram_n_41, A2 => gl_ram_ram_28(0), B1 => gl_ram_n_39, B2 => gl_ram_ram_27(0), ZN => gl_ram_n_82);
  gl_ram_g28807 : AOI22D0BWP7T port map(A1 => gl_ram_n_30, A2 => gl_ram_ram_89(0), B1 => gl_ram_n_29, B2 => gl_ram_ram_95(0), ZN => gl_ram_n_81);
  gl_ram_g28808 : AOI22D0BWP7T port map(A1 => gl_ram_n_41, A2 => gl_ram_ram_76(2), B1 => gl_ram_n_30, B2 => gl_ram_ram_73(2), ZN => gl_ram_n_80);
  gl_ram_g28809 : AOI22D0BWP7T port map(A1 => gl_ram_n_28, A2 => gl_ram_ram_82(2), B1 => gl_ram_n_31, B2 => gl_ram_ram_86(2), ZN => gl_ram_n_79);
  gl_ram_g28810 : AOI22D0BWP7T port map(A1 => gl_ram_n_30, A2 => gl_ram_ram_33(2), B1 => gl_ram_n_29, B2 => gl_ram_ram_39(2), ZN => gl_ram_n_78);
  gl_ram_g28811 : AOI22D0BWP7T port map(A1 => gl_ram_n_38, A2 => gl_ram_ram_80(2), B1 => gl_ram_n_29, B2 => gl_ram_ram_87(2), ZN => gl_ram_n_77);
  gl_ram_g28812 : AOI22D0BWP7T port map(A1 => gl_ram_n_41, A2 => gl_ram_ram_84(2), B1 => gl_ram_n_30, B2 => gl_ram_ram_81(2), ZN => gl_ram_n_76);
  gl_ram_g28813 : AOI22D0BWP7T port map(A1 => gl_ram_n_38, A2 => gl_ram_ram_40(0), B1 => gl_ram_n_29, B2 => gl_ram_ram_47(0), ZN => gl_ram_n_75);
  gl_ram_g28814 : AOI22D0BWP7T port map(A1 => gl_ram_n_28, A2 => gl_ram_ram_66(2), B1 => gl_ram_n_31, B2 => gl_ram_ram_70(2), ZN => gl_ram_n_74);
  gl_ram_g28815 : AOI22D0BWP7T port map(A1 => gl_ram_n_41, A2 => gl_ram_ram_44(0), B1 => gl_ram_n_30, B2 => gl_ram_ram_41(0), ZN => gl_ram_n_73);
  gl_ram_g28816 : AOI22D0BWP7T port map(A1 => gl_ram_n_28, A2 => gl_ram_ram_90(0), B1 => gl_ram_n_31, B2 => gl_ram_ram_94(0), ZN => gl_ram_n_72);
  gl_ram_g28817 : AOI22D0BWP7T port map(A1 => gl_ram_n_38, A2 => gl_ram_ram_64(2), B1 => gl_ram_n_29, B2 => gl_ram_ram_71(2), ZN => gl_ram_n_71);
  gl_ram_g28818 : AOI22D0BWP7T port map(A1 => gl_ram_n_40, A2 => gl_ram_ram_77(0), B1 => gl_ram_n_39, B2 => gl_ram_ram_75(0), ZN => gl_ram_n_70);
  gl_ram_g28819 : AOI22D0BWP7T port map(A1 => gl_ram_n_40, A2 => gl_ram_ram_61(2), B1 => gl_ram_n_39, B2 => gl_ram_ram_59(2), ZN => gl_ram_n_69);
  gl_ram_g28820 : AOI22D0BWP7T port map(A1 => gl_ram_n_30, A2 => gl_ram_ram_57(2), B1 => gl_ram_n_29, B2 => gl_ram_ram_63(2), ZN => gl_ram_n_68);
  gl_ram_g28821 : AOI22D0BWP7T port map(A1 => gl_ram_n_38, A2 => gl_ram_ram_72(0), B1 => gl_ram_n_41, B2 => gl_ram_ram_76(0), ZN => gl_ram_n_67);
  gl_ram_g28822 : AOI22D0BWP7T port map(A1 => gl_ram_n_28, A2 => gl_ram_ram_74(0), B1 => gl_ram_n_31, B2 => gl_ram_ram_78(0), ZN => gl_ram_n_66);
  gl_ram_g28823 : AOI22D0BWP7T port map(A1 => gl_ram_n_28, A2 => gl_ram_ram_58(2), B1 => gl_ram_n_31, B2 => gl_ram_ram_62(2), ZN => gl_ram_n_65);
  gl_ram_g28824 : AOI22D0BWP7T port map(A1 => gl_ram_n_38, A2 => gl_ram_ram_56(2), B1 => gl_ram_n_41, B2 => gl_ram_ram_60(2), ZN => gl_ram_n_64);
  gl_ram_g28825 : AOI22D0BWP7T port map(A1 => gl_ram_n_40, A2 => gl_ram_ram_13(2), B1 => gl_ram_n_39, B2 => gl_ram_ram_11(2), ZN => gl_ram_n_63);
  gl_ram_g28826 : AOI22D0BWP7T port map(A1 => gl_ram_n_30, A2 => gl_ram_ram_25(2), B1 => gl_ram_n_29, B2 => gl_ram_ram_31(2), ZN => gl_ram_n_62);
  gl_ram_g28827 : AOI22D0BWP7T port map(A1 => gl_ram_n_28, A2 => gl_ram_ram_74(1), B1 => gl_ram_n_31, B2 => gl_ram_ram_78(1), ZN => gl_ram_n_61);
  gl_ram_g28828 : HA1D0BWP7T port map(A => gl_ram_y_grid(1), B => gl_ram_y_grid(3), CO => gl_ram_n_56, S => gl_ram_n_57);
  gl_ram_g28829 : HA1D0BWP7T port map(A => gl_ram_x_grid(3), B => gl_ram_y_grid(0), CO => gl_ram_n_54, S => gl_ram_n_55);
  gl_ram_g28830 : IND2D1BWP7T port map(A1 => gl_ram_n_49, B1 => gl_ram_ram_position(5), ZN => gl_ram_n_60);
  gl_ram_g28831 : NR2XD0BWP7T port map(A1 => gl_ram_ram_position(5), A2 => gl_ram_n_49, ZN => gl_ram_n_59);
  gl_ram_g28832 : AN2D1BWP7T port map(A1 => gl_ram_n_32, A2 => gl_ram_n_20, Z => gl_ram_n_58);
  gl_ram_g28833 : INR2D1BWP7T port map(A1 => gl_ram_n_32, B1 => gl_ram_n_14, ZN => gl_ram_n_53);
  gl_ram_g28834 : AN2D1BWP7T port map(A1 => gl_ram_n_32, A2 => gl_ram_n_12, Z => gl_ram_n_52);
  gl_ram_g28835 : INR2D1BWP7T port map(A1 => gl_ram_n_32, B1 => gl_ram_n_13, ZN => gl_ram_n_51);
  gl_ram_g28836 : INVD1BWP7T port map(I => gl_ram_n_47, ZN => gl_ram_n_46);
  gl_ram_g28837 : INVD1BWP7T port map(I => gl_ram_n_43, ZN => gl_ram_n_42);
  gl_ram_g28838 : IND2D1BWP7T port map(A1 => gl_ram_n_7, B1 => gl_ram_ram_position(6), ZN => gl_ram_n_50);
  gl_ram_g28839 : INR2D1BWP7T port map(A1 => sig_logic_y(1), B1 => gl_ram_n_22, ZN => gl_ram_n_49);
  gl_ram_g28840 : NR2D1BWP7T port map(A1 => gl_ram_n_25, A2 => gl_ram_ram_position(4), ZN => gl_ram_n_48);
  gl_ram_g28841 : IND2D1BWP7T port map(A1 => gl_ram_n_21, B1 => gl_ram_ram_position(3), ZN => gl_ram_n_47);
  gl_ram_g28842 : AN2D1BWP7T port map(A1 => gl_ram_n_24, A2 => gl_ram_ram_position(4), Z => gl_ram_n_45);
  gl_ram_g28843 : AN2D1BWP7T port map(A1 => gl_ram_n_24, A2 => gl_ram_n_1, Z => gl_ram_n_44);
  gl_ram_g28844 : NR2XD0BWP7T port map(A1 => gl_ram_ram_position(3), A2 => gl_ram_n_21, ZN => gl_ram_n_43);
  gl_ram_g28845 : AN2D1BWP7T port map(A1 => gl_ram_n_20, A2 => gl_ram_ram_position(2), Z => gl_ram_n_41);
  gl_ram_g28846 : AN2D1BWP7T port map(A1 => gl_ram_n_12, A2 => gl_ram_ram_position(2), Z => gl_ram_n_40);
  gl_ram_g28847 : NR2D1BWP7T port map(A1 => gl_ram_n_14, A2 => gl_ram_ram_position(2), ZN => gl_ram_n_39);
  gl_ram_g28848 : AN2D1BWP7T port map(A1 => gl_ram_n_20, A2 => gl_ram_n_2, Z => gl_ram_n_38);
  gl_ram_g28849 : MAOI22D0BWP7T port map(A1 => gl_ram_n_4, A2 => gl_ram_x_grid(1), B1 => gl_ram_n_4, B2 => gl_ram_x_grid(1), ZN => gl_ram_n_27);
  gl_ram_g28850 : AOI21D0BWP7T port map(A1 => sig_logic_x(0), A2 => sig_logic_x(1), B => gl_ram_n_19, ZN => gl_ram_n_26);
  gl_ram_g28851 : NR2D1BWP7T port map(A1 => gl_ram_n_23, A2 => gl_ram_n_1, ZN => gl_ram_n_37);
  gl_ram_g28852 : NR2D1BWP7T port map(A1 => gl_ram_n_25, A2 => gl_ram_n_1, ZN => gl_ram_n_36);
  gl_ram_g28853 : NR2D1BWP7T port map(A1 => gl_ram_n_7, A2 => gl_ram_ram_position(6), ZN => gl_ram_n_35);
  gl_ram_g28854 : NR2D1BWP7T port map(A1 => gl_ram_n_15, A2 => gl_ram_ram_position(4), ZN => gl_ram_n_34);
  gl_ram_g28855 : NR2D1BWP7T port map(A1 => gl_ram_n_15, A2 => gl_ram_n_1, ZN => gl_ram_n_33);
  gl_ram_g28856 : NR2D1BWP7T port map(A1 => gl_ram_n_23, A2 => gl_ram_ram_position(4), ZN => gl_ram_n_32);
  gl_ram_g28857 : NR2D1BWP7T port map(A1 => gl_ram_n_13, A2 => gl_ram_n_2, ZN => gl_ram_n_31);
  gl_ram_g28858 : AN2D1BWP7T port map(A1 => gl_ram_n_12, A2 => gl_ram_n_2, Z => gl_ram_n_30);
  gl_ram_g28859 : NR2D1BWP7T port map(A1 => gl_ram_n_14, A2 => gl_ram_n_2, ZN => gl_ram_n_29);
  gl_ram_g28860 : NR2D1BWP7T port map(A1 => gl_ram_n_13, A2 => gl_ram_ram_position(2), ZN => gl_ram_n_28);
  gl_ram_g28861 : INVD0BWP7T port map(I => gl_ram_n_18, ZN => gl_ram_n_17);
  gl_ram_g28862 : CKND2D1BWP7T port map(A1 => gl_ram_ram_position(3), A2 => gl_ram_ram_position(5), ZN => gl_ram_n_25);
  gl_ram_g28863 : NR2D0BWP7T port map(A1 => gl_ram_ram_position(3), A2 => gl_ram_ram_position(5), ZN => gl_ram_n_24);
  gl_ram_g28864 : IND2D1BWP7T port map(A1 => gl_ram_ram_position(3), B1 => gl_ram_ram_position(5), ZN => gl_ram_n_23);
  gl_ram_g28865 : ND2D1BWP7T port map(A1 => sig_logic_y(3), A2 => sig_logic_y(2), ZN => gl_ram_n_22);
  gl_ram_g28866 : INR2D1BWP7T port map(A1 => gl_ram_x_grid(1), B1 => gl_ram_n_4, ZN => gl_ram_n_16);
  gl_ram_g28867 : NR2XD0BWP7T port map(A1 => sig_logic_y(3), A2 => sig_logic_y(2), ZN => gl_ram_n_21);
  gl_ram_g28868 : NR2D0BWP7T port map(A1 => gl_ram_ram_position(0), A2 => gl_ram_ram_position(1), ZN => gl_ram_n_20);
  gl_ram_g28869 : NR2XD0BWP7T port map(A1 => sig_logic_x(0), A2 => sig_logic_x(1), ZN => gl_ram_n_19);
  gl_ram_g28870 : NR2D1BWP7T port map(A1 => sig_middelsteknop, A2 => gl_ram_ram_position(4), ZN => gl_ram_n_18);
  gl_ram_g28871 : IND2D1BWP7T port map(A1 => gl_ram_ram_position(5), B1 => gl_ram_ram_position(3), ZN => gl_ram_n_15);
  gl_ram_g28872 : ND2D1BWP7T port map(A1 => gl_ram_ram_position(1), A2 => gl_ram_ram_position(0), ZN => gl_ram_n_14);
  gl_ram_g28873 : ND2D1BWP7T port map(A1 => gl_ram_n_3, A2 => gl_ram_ram_position(1), ZN => gl_ram_n_13);
  gl_ram_g28874 : NR2D1BWP7T port map(A1 => gl_ram_n_3, A2 => gl_ram_ram_position(1), ZN => gl_ram_n_12);
  gl_ram_g28875 : NR2XD0BWP7T port map(A1 => gl_ram_ram_position(4), A2 => gl_ram_ram_position(0), ZN => gl_ram_n_11);
  gl_ram_g28876 : ND2D1BWP7T port map(A1 => gl_ram_ram_position(4), A2 => gl_ram_ram_position(0), ZN => gl_ram_n_10);
  gl_ram_g28877 : NR2XD0BWP7T port map(A1 => gl_ram_n_1, A2 => gl_ram_ram_position(0), ZN => gl_ram_n_9);
  gl_ram_g28878 : ND2D1BWP7T port map(A1 => gl_ram_n_1, A2 => gl_ram_ram_position(0), ZN => gl_ram_n_8);
  gl_ram_g28879 : CKAN2D1BWP7T port map(A1 => gl_sig_countdown_aan, A2 => sig_draw, Z => gl_ram_n_7);
  gl_ram_g28884 : INVD1BWP7T port map(I => sig_middelsteknop, ZN => gl_ram_n_6);
  gl_ram_g28885 : CKND1BWP7T port map(I => sig_logic_x(2), ZN => gl_ram_n_5);
  gl_ram_ram_position_reg_0 : DFD1BWP7T port map(CP => clk, D => gl_ram_n_457, Q => gl_ram_ram_position(0), QN => gl_ram_n_3);
  gl_ram_ram_position_reg_2 : DFD1BWP7T port map(CP => clk, D => gl_ram_n_454, Q => gl_ram_ram_position(2), QN => gl_ram_n_2);
  gl_ram_ram_position_reg_4 : DFD0BWP7T port map(CP => clk, D => gl_ram_n_468, Q => gl_ram_ram_position(4), QN => gl_ram_n_1);
  gl_ram_y_grid_reg_0 : DFD1BWP7T port map(CP => clk, D => gl_ram_n_461, Q => gl_ram_y_grid(0), QN => gl_ram_n_4);
  gl_ram_g14056 : IND2D1BWP7T port map(A1 => n_0, B1 => gl_ram_n_6, ZN => gl_ram_n_0);
  ml_g3 : BUFFD4BWP7T port map(I => ml_mouseX(1), Z => led8);
  ml_g1 : BUFFD4BWP7T port map(I => ml_buttons_mouse(4), Z => led5);
  ml_g2 : BUFFD4BWP7T port map(I => ml_buttons_mouse(1), Z => led0);
  ml_ms_g701 : BUFFD4BWP7T port map(I => ml_ms_n_82, Z => led6);
  ml_ms_g700 : BUFFD4BWP7T port map(I => ml_ms_n_78, Z => led9);
  ml_ms_g759 : OR2D4BWP7T port map(A1 => ml_ms_n_62, A2 => ml_ms_n_63, Z => clk15k_switch);
  ml_ms_g760 : INR2XD0BWP7T port map(A1 => ml_ms_sfsm_n_383, B1 => ml_ms_muxFSM, ZN => ml_ms_n_63);
  ml_ms_g762 : NR2XD0BWP7T port map(A1 => ml_ms_n_61, A2 => ml_ms_sfsm_state(0), ZN => ml_ms_n_62);
  ml_ms_g763 : CKAN2D1BWP7T port map(A1 => ml_ms_sfsm_state(1), A2 => ml_ms_sfsm_state(0), Z => ml_ms_sfsm_n_383);
  ml_ms_g765 : IND2D1BWP7T port map(A1 => ml_ms_sfsm_state(1), B1 => ml_ms_muxFSM, ZN => ml_ms_n_61);
  ml_ms_g2 : INR2D1BWP7T port map(A1 => ml_ms_n_61, B1 => ml_ms_sfsm_state(0), ZN => ml_ms_cntReset25M_send);
  ml_ms_sfsm_state_reg_0 : DFQD1BWP7T port map(CP => clk, D => ml_ms_n_58, Q => ml_ms_sfsm_state(0));
  ml_ms_sr_new_new_data_reg_0 : DFQD1BWP7T port map(CP => clk, D => ml_ms_n_30, Q => ml_ms_sr_new_new_data(0));
  ml_ms_sr_new_new_data_reg_1 : DFQD1BWP7T port map(CP => clk, D => ml_ms_n_20, Q => ml_ms_sr_new_new_data(1));
  ml_ms_sr_new_new_data_reg_2 : DFQD1BWP7T port map(CP => clk, D => ml_ms_n_19, Q => ml_ms_sr_new_new_data(2));
  ml_ms_sr_new_new_data_reg_3 : DFQD1BWP7T port map(CP => clk, D => ml_ms_n_26, Q => ml_ms_sr_new_new_data(3));
  ml_ms_sr_new_new_data_reg_4 : DFQD1BWP7T port map(CP => clk, D => ml_ms_n_25, Q => ml_ms_sr_new_new_data(4));
  ml_ms_sr_new_new_data_reg_5 : DFQD1BWP7T port map(CP => clk, D => ml_ms_n_34, Q => ml_ms_sr_new_new_data(5));
  ml_ms_sr_new_new_data_reg_6 : DFQD1BWP7T port map(CP => clk, D => ml_ms_n_24, Q => ml_ms_sr_new_new_data(6));
  ml_ms_sr_new_new_data_reg_7 : DFQD1BWP7T port map(CP => clk, D => ml_ms_n_32, Q => ml_ms_sr_new_new_data(7));
  ml_ms_sr_new_new_data_reg_8 : DFQD1BWP7T port map(CP => clk, D => ml_ms_n_31, Q => ml_ms_muxReg);
  ml_ms_g1851 : MOAI22D0BWP7T port map(A1 => ml_ms_n_45, A2 => ml_ms_n_10, B1 => ml_ms_n_59, B2 => ml_ms_mux_select, ZN => ml_ms_n_60);
  ml_ms_g1854 : OAI211D1BWP7T port map(A1 => ml_ms_n_8, A2 => ml_ms_n_47, B => ml_ms_n_52, C => ml_ms_n_55, ZN => ml_ms_n_59);
  ml_ms_g1855 : OAI211D1BWP7T port map(A1 => ml_ms_n_49, A2 => ml_ms_n_53, B => ml_ms_n_52, C => ml_ms_n_56, ZN => ml_ms_n_58);
  ml_ms_g1856 : OAI221D0BWP7T port map(A1 => ml_ms_n_53, A2 => ml_ms_n_50, B1 => ml_ms_n_0, B2 => ml_ms_n_8, C => ml_ms_n_51, ZN => ml_ms_n_57);
  ml_ms_g1858 : OAI21D0BWP7T port map(A1 => ml_ms_n_47, A2 => ml_ms_n_14, B => ml_ms_n_7, ZN => ml_ms_n_56);
  ml_ms_g1859 : IND3D1BWP7T port map(A1 => ml_ms_n_10, B1 => ml_ms_muxFSM, B2 => ml_ms_n_50, ZN => ml_ms_n_55);
  ml_ms_g1860 : MOAI22D0BWP7T port map(A1 => ml_ms_n_48, A2 => ml_ms_n_16, B1 => ml_ms_n_46, B2 => ml_ms_muxFSM, ZN => ml_ms_n_54);
  ml_ms_g1861 : IND3D1BWP7T port map(A1 => ml_ms_n_10, B1 => ml_ms_muxFSM, B2 => ml_ms_n_45, ZN => ml_ms_n_53);
  ml_ms_g1862 : IND3D1BWP7T port map(A1 => ml_ms_n_40, B1 => ml_ms_n_45, B2 => ml_ms_n_48, ZN => ml_ms_n_51);
  ml_ms_g1863 : IND3D1BWP7T port map(A1 => ml_ms_n_16, B1 => ml_ms_n_37, B2 => ml_ms_n_48, ZN => ml_ms_n_52);
  ml_ms_g1864 : INVD0BWP7T port map(I => ml_ms_n_50, ZN => ml_ms_n_49);
  ml_ms_g1865 : IAO21D0BWP7T port map(A1 => ml_ms_n_43, A2 => ml_ms_n_11, B => ml_ms_count25M(12), ZN => ml_ms_n_50);
  ml_ms_g1866 : IOA21D1BWP7T port map(A1 => ml_ms_n_42, A2 => ml_ms_n_18, B => ml_ms_sfsm_state(1), ZN => ml_ms_n_48);
  ml_ms_g1867 : AOI21D0BWP7T port map(A1 => ml_ms_n_44, A2 => ml_ms_sfsm_state(0), B => ml_ms_reset_send, ZN => ml_ms_n_46);
  ml_ms_g1868 : AOI211XD0BWP7T port map(A1 => ml_ms_sfsm_state(1), A2 => ml_ms_Clk15k_buffered, B => ml_ms_n_41, C => ml_ms_n_1, ZN => ml_ms_n_47);
  ml_ms_g1869 : ND2D1BWP7T port map(A1 => ml_ms_n_44, A2 => ml_ms_muxFSM, ZN => ml_ms_n_45);
  ml_ms_g1870 : NR2XD0BWP7T port map(A1 => ml_ms_n_38, A2 => ml_ms_count25M(9), ZN => ml_ms_n_43);
  ml_ms_g1871 : OA31D1BWP7T port map(A1 => ml_ms_count25M(11), A2 => ml_ms_count25M(10), A3 => ml_ms_n_33, B => ml_ms_sfsm_state(1), Z => ml_ms_n_44);
  ml_ms_g1872 : OAI211D1BWP7T port map(A1 => ml_ms_n_17, A2 => ml_ms_n_36, B => ml_ms_count25M(11), C => ml_ms_count25M(9), ZN => ml_ms_n_42);
  ml_ms_g1873 : NR2D1BWP7T port map(A1 => ml_ms_n_39, A2 => ml_ms_sfsm_state(1), ZN => ml_ms_n_41);
  ml_ms_g1874 : OA22D0BWP7T port map(A1 => ml_ms_n_16, A2 => ml_ms_n_37, B1 => ml_ms_n_0, B2 => ml_ms_n_10, Z => ml_ms_n_40);
  ml_ms_g1875 : AOI21D0BWP7T port map(A1 => ml_ms_n_35, A2 => ml_ms_n_15, B => ml_ms_n_18, ZN => ml_ms_n_39);
  ml_ms_g1876 : AO211D0BWP7T port map(A1 => ml_ms_n_27, A2 => ml_ms_count25M(8), B => ml_ms_n_29, C => ml_ms_n_17, Z => ml_ms_n_38);
  ml_ms_g1881 : ND4D0BWP7T port map(A1 => ml_ms_n_12, A2 => ml_ms_count25M(8), A3 => ml_ms_count25M(9), A4 => ml_ms_count25M(12), ZN => ml_ms_n_37);
  ml_ms_g1882 : AN2D0BWP7T port map(A1 => ml_ms_n_29, A2 => ml_ms_count25M(3), Z => ml_ms_n_36);
  ml_ms_g1888 : OAI211D1BWP7T port map(A1 => ml_ms_count25M(3), A2 => ml_ms_n_3, B => ml_ms_n_5, C => ml_ms_count25M(5), ZN => ml_ms_n_35);
  ml_ms_g1889 : ND2D1BWP7T port map(A1 => ml_ms_n_28, A2 => ml_ms_n_22, ZN => ml_ms_n_34);
  ml_ms_g1890 : OAI21D0BWP7T port map(A1 => ml_ms_n_13, A2 => ml_ms_n_6, B => ml_ms_n_15, ZN => ml_ms_n_33);
  ml_ms_g1891 : ND2D1BWP7T port map(A1 => ml_ms_n_28, A2 => ml_ms_n_23, ZN => ml_ms_n_32);
  ml_ms_g1892 : ND2D1BWP7T port map(A1 => ml_ms_n_28, A2 => ml_ms_n_21, ZN => ml_ms_n_31);
  ml_ms_g1893 : IOA21D1BWP7T port map(A1 => ml_ms_n_4, A2 => ml_ms_sr_new_new_data(0), B => ml_ms_n_28, ZN => ml_ms_n_30);
  ml_ms_g1894 : AN4D0BWP7T port map(A1 => ml_ms_count25M(3), A2 => ml_ms_count25M(2), A3 => ml_ms_count25M(7), A4 => ml_ms_count25M(5), Z => ml_ms_n_27);
  ml_ms_g1895 : AO22D0BWP7T port map(A1 => ml_ms_n_4, A2 => ml_ms_sr_new_new_data(3), B1 => ml_ms_sr_new_new_data(2), B2 => ml_ms_n_9, Z => ml_ms_n_26);
  ml_ms_g1896 : AO22D0BWP7T port map(A1 => ml_ms_n_4, A2 => ml_ms_sr_new_new_data(4), B1 => ml_ms_sr_new_new_data(3), B2 => ml_ms_n_9, Z => ml_ms_n_25);
  ml_ms_g1897 : AN4D0BWP7T port map(A1 => ml_ms_count25M(4), A2 => ml_ms_count25M(8), A3 => ml_ms_count25M(7), A4 => ml_ms_count25M(5), Z => ml_ms_n_29);
  ml_ms_g1898 : OAI211D1BWP7T port map(A1 => ml_ms_muxFSM, A2 => ml_ms_sfsm_n_383, B => ml_ms_actBit, C => ml_ms_n_2, ZN => ml_ms_n_28);
  ml_ms_g1899 : AO22D0BWP7T port map(A1 => ml_ms_n_4, A2 => ml_ms_sr_new_new_data(6), B1 => ml_ms_sr_new_new_data(5), B2 => ml_ms_n_9, Z => ml_ms_n_24);
  ml_ms_g1900 : AOI22D0BWP7T port map(A1 => ml_ms_n_4, A2 => ml_ms_sr_new_new_data(7), B1 => ml_ms_n_9, B2 => ml_ms_sr_new_new_data(6), ZN => ml_ms_n_23);
  ml_ms_g1901 : AOI22D0BWP7T port map(A1 => ml_ms_n_4, A2 => ml_ms_sr_new_new_data(5), B1 => ml_ms_n_9, B2 => ml_ms_sr_new_new_data(4), ZN => ml_ms_n_22);
  ml_ms_g1902 : AOI22D0BWP7T port map(A1 => ml_ms_n_4, A2 => ml_ms_muxReg, B1 => ml_ms_n_9, B2 => ml_ms_sr_new_new_data(7), ZN => ml_ms_n_21);
  ml_ms_g1903 : AO22D0BWP7T port map(A1 => ml_ms_n_4, A2 => ml_ms_sr_new_new_data(1), B1 => ml_ms_sr_new_new_data(0), B2 => ml_ms_n_9, Z => ml_ms_n_20);
  ml_ms_g1904 : AO22D0BWP7T port map(A1 => ml_ms_n_4, A2 => ml_ms_sr_new_new_data(2), B1 => ml_ms_sr_new_new_data(1), B2 => ml_ms_n_9, Z => ml_ms_n_19);
  ml_ms_g1905 : INR2D1BWP7T port map(A1 => ml_ms_n_11, B1 => ml_ms_count25M(12), ZN => ml_ms_n_18);
  ml_ms_g1906 : INR2D1BWP7T port map(A1 => ml_ms_count25M(8), B1 => ml_ms_n_6, ZN => ml_ms_n_17);
  ml_ms_g1907 : OR2D1BWP7T port map(A1 => ml_ms_n_10, A2 => ml_ms_muxFSM, Z => ml_ms_n_16);
  ml_ms_g1908 : AOI21D0BWP7T port map(A1 => ml_ms_n_0, A2 => ml_ms_mux_select, B => ml_ms_muxFSM, ZN => ml_ms_n_14);
  ml_ms_g1909 : NR3D0BWP7T port map(A1 => ml_ms_count25M(3), A2 => ml_ms_count25M(4), A3 => ml_ms_count25M(5), ZN => ml_ms_n_13);
  ml_ms_g1910 : IAO21D0BWP7T port map(A1 => ml_ms_count25M(7), A2 => ml_ms_count25M(6), B => ml_ms_n_11, ZN => ml_ms_n_12);
  ml_ms_g1911 : NR3D0BWP7T port map(A1 => ml_ms_count25M(8), A2 => ml_ms_count25M(12), A3 => ml_ms_count25M(9), ZN => ml_ms_n_15);
  ml_ms_g1912 : ND2D1BWP7T port map(A1 => ml_ms_count25M(10), A2 => ml_ms_count25M(11), ZN => ml_ms_n_11);
  ml_ms_g1913 : IND2D1BWP7T port map(A1 => ml_ms_reset_send, B1 => ml_ms_sfsm_state(0), ZN => ml_ms_n_10);
  ml_ms_g1914 : AN2D1BWP7T port map(A1 => ml_ms_output_edgedet, A2 => ml_ms_mux_select, Z => ml_ms_n_9);
  ml_ms_g1915 : INVD1BWP7T port map(I => ml_ms_n_7, ZN => ml_ms_n_8);
  ml_ms_g1916 : INVD0BWP7T port map(I => ml_ms_n_6, ZN => ml_ms_n_5);
  ml_ms_g1917 : OR2D1BWP7T port map(A1 => ml_ms_count25M(4), A2 => ml_ms_count25M(2), Z => ml_ms_n_3);
  ml_ms_g1918 : NR2XD0BWP7T port map(A1 => ml_ms_reset_send, A2 => ml_ms_sfsm_state(0), ZN => ml_ms_n_7);
  ml_ms_g1919 : CKND2D1BWP7T port map(A1 => ml_ms_count25M(7), A2 => ml_ms_count25M(6), ZN => ml_ms_n_6);
  ml_ms_g1920 : NR2XD0BWP7T port map(A1 => ml_ms_output_edgedet, A2 => ml_ms_n_2, ZN => ml_ms_n_4);
  ml_ms_sfsm_state_reg_1 : DFD1BWP7T port map(CP => clk, D => ml_ms_n_57, Q => ml_ms_sfsm_state(1), QN => ml_ms_n_0);
  ml_ms_sfsm_state_reg_3 : DFD1BWP7T port map(CP => clk, D => ml_ms_n_60, Q => ml_ms_mux_select, QN => ml_ms_n_2);
  ml_ms_sfsm_state_reg_2 : DFD1BWP7T port map(CP => clk, D => ml_ms_n_54, Q => ml_ms_muxFSM, QN => ml_ms_n_1);
  ml_ms_mfsm_g2695 : MOAI22D0BWP7T port map(A1 => ml_ms_mfsm_n_75, A2 => ml_ms_data_sr_11bit(4), B1 => ml_ms_mfsm_n_74, B2 => ml_ms_data_sr_11bit(4), ZN => ml_ms_mouse_x(2));
  ml_ms_mfsm_g2696 : MOAI22D0BWP7T port map(A1 => ml_ms_mfsm_n_75, A2 => ml_ms_data_sr_11bit(5), B1 => ml_ms_mfsm_n_74, B2 => ml_ms_data_sr_11bit(5), ZN => ml_ms_mouse_x(1));
  ml_ms_mfsm_g2697 : MOAI22D0BWP7T port map(A1 => ml_ms_mfsm_n_75, A2 => ml_ms_data_sr_11bit(6), B1 => ml_ms_mfsm_n_74, B2 => ml_ms_data_sr_11bit(6), ZN => ml_ms_mouse_x(0));
  ml_ms_mfsm_g2698 : MOAI22D0BWP7T port map(A1 => ml_ms_mfsm_n_73, A2 => ml_ms_data_sr_11bit(4), B1 => ml_ms_mfsm_n_72, B2 => ml_ms_data_sr_11bit(4), ZN => ml_ms_mouse_y(2));
  ml_ms_mfsm_g2699 : MOAI22D0BWP7T port map(A1 => ml_ms_mfsm_n_73, A2 => ml_ms_data_sr_11bit(5), B1 => ml_ms_mfsm_n_72, B2 => ml_ms_data_sr_11bit(5), ZN => ml_ms_mouse_y(1));
  ml_ms_mfsm_g2700 : MOAI22D0BWP7T port map(A1 => ml_ms_mfsm_n_73, A2 => ml_ms_data_sr_11bit(6), B1 => ml_ms_mfsm_n_72, B2 => ml_ms_data_sr_11bit(6), ZN => ml_ms_mouse_y(0));
  ml_ms_mfsm_g2701 : AO21D0BWP7T port map(A1 => ml_ms_mfsm_state(3), A2 => ml_ms_mfsm_n_69, B => ml_ms_mux_select_main, Z => ml_ms_timerReset);
  ml_ms_mfsm_g2702 : ND2D1BWP7T port map(A1 => ml_ms_mfsm_n_70, A2 => ml_ms_n_82, ZN => ml_ms_mfsm_n_75);
  ml_ms_mfsm_g2703 : NR2D1BWP7T port map(A1 => ml_ms_n_82, A2 => ml_ms_mfsm_n_71, ZN => ml_ms_mfsm_n_74);
  ml_ms_mfsm_g2704 : IND3D1BWP7T port map(A1 => ml_ms_mfsm_n_60, B1 => ml_ms_mfsm_n_67, B2 => ml_buttons_mouse(1), ZN => ml_ms_mfsm_n_73);
  ml_ms_mfsm_g2705 : NR3D0BWP7T port map(A1 => ml_ms_mfsm_n_60, A2 => ml_buttons_mouse(1), A3 => ml_ms_mfsm_n_68, ZN => ml_ms_mfsm_n_72);
  ml_ms_mfsm_g2706 : CKND1BWP7T port map(I => ml_ms_mfsm_n_70, ZN => ml_ms_mfsm_n_71);
  ml_ms_mfsm_g2707 : NR2XD0BWP7T port map(A1 => ml_ms_mfsm_n_58, A2 => ml_ms_mfsm_n_68, ZN => ml_ms_mfsm_n_70);
  ml_ms_mfsm_g2708 : OAI21D0BWP7T port map(A1 => ml_ms_mfsm_n_45, A2 => ml_ms_mfsm_n_66, B => ml_ms_mfsm_n_52, ZN => ml_ms_mfsm_n_69);
  ml_ms_mfsm_g2709 : INVD1BWP7T port map(I => ml_ms_mfsm_n_67, ZN => ml_ms_mfsm_n_68);
  ml_ms_mfsm_g2710 : NR2XD0BWP7T port map(A1 => ml_ms_mfsm_n_0, A2 => ml_ms_mfsm_n_66, ZN => ml_ms_mfsm_n_67);
  ml_ms_mfsm_g2711 : OAI31D0BWP7T port map(A1 => ml_ms_timer_count(20), A2 => ml_ms_timer_count(19), A3 => ml_ms_mfsm_n_65, B => ml_ms_timer_count(21), ZN => ml_ms_mfsm_n_66);
  ml_ms_mfsm_g2712 : AN3D0BWP7T port map(A1 => ml_ms_mfsm_n_64, A2 => ml_ms_timer_count(18), A3 => ml_ms_timer_count(17), Z => ml_ms_mfsm_n_65);
  ml_ms_mfsm_g2713 : OR4D0BWP7T port map(A1 => ml_ms_timer_count(16), A2 => ml_ms_timer_count(14), A3 => ml_ms_timer_count(15), A4 => ml_ms_mfsm_n_63, Z => ml_ms_mfsm_n_64);
  ml_ms_mfsm_g2714 : OA31D0BWP7T port map(A1 => ml_ms_timer_count(12), A2 => ml_ms_timer_count(11), A3 => ml_ms_mfsm_n_62, B => ml_ms_timer_count(13), Z => ml_ms_mfsm_n_63);
  ml_ms_mfsm_g2715 : AN2D0BWP7T port map(A1 => ml_ms_btnflipfloprst, A2 => ml_ms_data_sr_11bit(8), Z => ml_ms_btns(4));
  ml_ms_mfsm_g2716 : AN2D0BWP7T port map(A1 => ml_ms_btnflipfloprst, A2 => ml_ms_data_sr_11bit(7), Z => ml_ms_btns(3));
  ml_ms_mfsm_g2717 : AN2D0BWP7T port map(A1 => ml_ms_btnflipfloprst, A2 => ml_ms_data_sr_11bit(9), Z => ml_ms_btns(2));
  ml_ms_mfsm_g2718 : AN2D0BWP7T port map(A1 => ml_ms_btnflipfloprst, A2 => ml_ms_data_sr_11bit(4), Z => ml_ms_btns(1));
  ml_ms_mfsm_g2719 : AN2D0BWP7T port map(A1 => ml_ms_btnflipfloprst, A2 => ml_ms_data_sr_11bit(5), Z => ml_ms_btns(0));
  ml_ms_mfsm_g2720 : ND3D0BWP7T port map(A1 => ml_ms_mfsm_n_56, A2 => ml_ms_mfsm_n_59, A3 => ml_ms_mfsm_state(1), ZN => ml_ms_cntReset25M_main);
  ml_ms_mfsm_g2721 : OAI211D1BWP7T port map(A1 => ml_ms_mfsm_state(0), A2 => ml_ms_mfsm_n_54, B => ml_ms_mfsm_n_61, C => ml_ms_mfsm_n_53, ZN => ml_ms_cntReset15K);
  ml_ms_mfsm_g2722 : MOAI22D0BWP7T port map(A1 => ml_ms_mfsm_n_50, A2 => ml_ms_mfsm_n_47, B1 => ml_ms_mfsm_n_57, B2 => ml_ms_mfsm_state(4), ZN => ml_ms_btnflipfloprst);
  ml_ms_mfsm_g2723 : NR2XD0BWP7T port map(A1 => ml_ms_mfsm_n_60, A2 => ml_ms_mfsm_n_0, ZN => ml_ms_yflipfloprst);
  ml_ms_mfsm_g2724 : OA21D0BWP7T port map(A1 => ml_ms_mfsm_n_51, A2 => ml_ms_timer_count(9), B => ml_ms_timer_count(10), Z => ml_ms_mfsm_n_62);
  ml_ms_mfsm_g2725 : AOI22D0BWP7T port map(A1 => ml_ms_mfsm_n_54, A2 => ml_ms_mfsm_n_48, B1 => ml_ms_mfsm_state(4), B2 => ml_ms_mfsm_state(3), ZN => ml_ms_mfsm_n_61);
  ml_ms_mfsm_g2726 : NR2XD0BWP7T port map(A1 => ml_ms_mfsm_n_52, A2 => ml_ms_mfsm_n_0, ZN => ml_ms_xflipfloprst);
  ml_ms_mfsm_g2727 : ND2D1BWP7T port map(A1 => ml_ms_mfsm_n_55, A2 => ml_ms_mfsm_state(0), ZN => ml_ms_reset_send);
  ml_ms_mfsm_g2729 : ND2D1BWP7T port map(A1 => ml_ms_mfsm_n_53, A2 => ml_ms_mfsm_n_54, ZN => ml_ms_mux_select_main);
  ml_ms_mfsm_g2730 : AOI32D1BWP7T port map(A1 => ml_ms_mfsm_n_43, A2 => ml_ms_mfsm_n_0, A3 => ml_ms_mfsm_state(2), B1 => ml_ms_mfsm_n_1, B2 => ml_ms_mfsm_state(3), ZN => ml_ms_mfsm_n_59);
  ml_ms_mfsm_g2731 : OA21D0BWP7T port map(A1 => ml_ms_mfsm_n_45, A2 => ml_ms_mfsm_n_1, B => ml_ms_mfsm_n_52, Z => ml_ms_mfsm_n_58);
  ml_ms_mfsm_g2732 : NR3D0BWP7T port map(A1 => ml_ms_mfsm_n_45, A2 => ml_ms_mfsm_state(3), A3 => ml_ms_mfsm_state(2), ZN => ml_ms_mfsm_n_57);
  ml_ms_mfsm_g2733 : MAOI22D0BWP7T port map(A1 => ml_ms_mfsm_n_49, A2 => ml_ms_mfsm_state(0), B1 => ml_ms_mfsm_n_49, B2 => ml_ms_mfsm_state(0), ZN => ml_ms_mfsm_n_56);
  ml_ms_mfsm_g2734 : AOI22D0BWP7T port map(A1 => ml_ms_mfsm_n_46, A2 => ml_ms_mfsm_state(3), B1 => ml_ms_mfsm_n_48, B2 => ml_ms_mfsm_state(2), ZN => ml_ms_mfsm_n_60);
  ml_ms_mfsm_g2736 : AN2D1BWP7T port map(A1 => ml_ms_mfsm_n_148, A2 => ml_ms_mfsm_state(4), Z => ml_handshake_mouse_out);
  ml_ms_mfsm_g2737 : NR2XD0BWP7T port map(A1 => ml_ms_mfsm_n_49, A2 => ml_ms_mfsm_state(1), ZN => ml_ms_mfsm_n_55);
  ml_ms_mfsm_g2738 : ND2D1BWP7T port map(A1 => ml_ms_mfsm_n_50, A2 => ml_ms_mfsm_n_0, ZN => ml_ms_mfsm_n_54);
  ml_ms_mfsm_g2739 : OA211D0BWP7T port map(A1 => ml_ms_timer_count(5), A2 => ml_ms_timer_count(6), B => ml_ms_timer_count(8), C => ml_ms_timer_count(7), Z => ml_ms_mfsm_n_51);
  ml_ms_mfsm_g2740 : ND2D1BWP7T port map(A1 => ml_ms_mfsm_n_46, A2 => ml_ms_mfsm_n_0, ZN => ml_ms_mfsm_n_53);
  ml_ms_mfsm_g2741 : ND2D1BWP7T port map(A1 => ml_ms_mfsm_n_48, A2 => ml_ms_mfsm_n_1, ZN => ml_ms_mfsm_n_52);
  ml_ms_mfsm_g2742 : ND2D1BWP7T port map(A1 => ml_ms_mfsm_state(3), A2 => ml_ms_mfsm_state(2), ZN => ml_ms_mfsm_n_50);
  ml_ms_mfsm_g2743 : INR2D1BWP7T port map(A1 => ml_ms_mfsm_state(0), B1 => ml_ms_mfsm_n_43, ZN => ml_ms_mfsm_n_148);
  ml_ms_mfsm_g2744 : INVD0BWP7T port map(I => ml_ms_mfsm_n_47, ZN => ml_ms_mfsm_n_48);
  ml_ms_mfsm_g2745 : INVD1BWP7T port map(I => ml_ms_mfsm_n_46, ZN => ml_ms_mfsm_n_45);
  ml_ms_mfsm_g2746 : ND2D1BWP7T port map(A1 => ml_ms_mfsm_n_1, A2 => ml_ms_mfsm_n_0, ZN => ml_ms_mfsm_n_49);
  ml_ms_mfsm_g2747 : ND2D1BWP7T port map(A1 => ml_ms_mfsm_state(0), A2 => ml_ms_mfsm_state(1), ZN => ml_ms_mfsm_n_47);
  ml_ms_mfsm_g2748 : NR2XD0BWP7T port map(A1 => ml_ms_mfsm_state(0), A2 => ml_ms_mfsm_state(1), ZN => ml_ms_mfsm_n_46);
  ml_ms_mfsm_g2 : CKAN2D1BWP7T port map(A1 => ml_ms_mfsm_n_148, A2 => ml_ms_mfsm_n_55, Z => ml_ms_actBit);
  ml_ms_mfsm_state_reg_0 : DFQD1BWP7T port map(CP => clk, D => ml_ms_mfsm_n_40, Q => ml_ms_mfsm_state(0));
  ml_ms_mfsm_state_reg_1 : DFQD1BWP7T port map(CP => clk, D => ml_ms_mfsm_n_41, Q => ml_ms_mfsm_state(1));
  ml_ms_mfsm_g2795 : OAI21D0BWP7T port map(A1 => ml_ms_mfsm_n_27, A2 => ml_ms_mfsm_state(1), B => ml_ms_mfsm_n_39, ZN => ml_ms_mfsm_n_41);
  ml_ms_mfsm_g2796 : AO33D0BWP7T port map(A1 => ml_ms_mfsm_n_38, A2 => ml_ms_mfsm_n_13, A3 => ml_ms_mfsm_state(1), B1 => ml_ms_mfsm_n_33, B2 => ml_ms_mfsm_n_12, B3 => ml_ms_mfsm_n_5, Z => ml_ms_mfsm_n_40);
  ml_ms_mfsm_g2797 : ND4D0BWP7T port map(A1 => ml_ms_mfsm_n_36, A2 => ml_ms_mfsm_n_22, A3 => ml_ms_mfsm_n_11, A4 => ml_ms_mfsm_state(1), ZN => ml_ms_mfsm_n_39);
  ml_ms_mfsm_g2799 : AOI21D0BWP7T port map(A1 => ml_ms_mfsm_n_30, A2 => ml_ms_mfsm_n_3, B => ml_ms_mfsm_n_37, ZN => ml_ms_mfsm_n_38);
  ml_ms_mfsm_g2800 : AOI21D0BWP7T port map(A1 => ml_ms_mfsm_n_35, A2 => ml_ms_mfsm_n_22, B => ml_ms_mfsm_state(4), ZN => ml_ms_mfsm_n_37);
  ml_ms_mfsm_g2801 : AOI32D1BWP7T port map(A1 => ml_ms_mfsm_n_32, A2 => ml_ms_mfsm_state(4), A3 => ml_ms_mfsm_state(3), B1 => ml_ms_mfsm_n_25, B2 => ml_ms_mfsm_state(2), ZN => ml_ms_mfsm_n_36);
  ml_ms_mfsm_g2802 : OAI211D1BWP7T port map(A1 => ml_ms_mfsm_state(0), A2 => ml_ms_mfsm_n_30, B => ml_ms_mfsm_state(2), C => ml_ms_mfsm_state(3), ZN => ml_ms_mfsm_n_35);
  ml_ms_mfsm_g2803 : AOI22D0BWP7T port map(A1 => ml_ms_mfsm_n_31, A2 => ml_ms_mfsm_state(2), B1 => ml_ms_mfsm_n_28, B2 => ml_ms_mfsm_n_1, ZN => ml_ms_mfsm_n_34);
  ml_ms_mfsm_g2805 : OAI22D0BWP7T port map(A1 => ml_ms_mfsm_n_29, A2 => ml_ms_mfsm_state(2), B1 => ml_ms_mfsm_n_21, B2 => ml_ms_mfsm_n_1, ZN => ml_ms_mfsm_n_33);
  ml_ms_mfsm_g2806 : OAI22D0BWP7T port map(A1 => ml_ms_mfsm_n_30, A2 => ml_ms_mfsm_n_1, B1 => ml_ms_mfsm_state(0), B2 => ml_ms_mfsm_state(2), ZN => ml_ms_mfsm_n_32);
  ml_ms_mfsm_g2807 : IOA21D1BWP7T port map(A1 => ml_ms_mfsm_n_25, A2 => ml_ms_mfsm_n_0, B => ml_ms_mfsm_n_13, ZN => ml_ms_mfsm_n_31);
  ml_ms_mfsm_g2808 : AN2D0BWP7T port map(A1 => ml_ms_mfsm_n_25, A2 => ml_ms_mfsm_state(4), Z => ml_ms_mfsm_n_29);
  ml_ms_mfsm_g2809 : INR2D1BWP7T port map(A1 => ml_ms_mfsm_n_23, B1 => ml_ms_count25M(12), ZN => ml_ms_mfsm_n_30);
  ml_ms_mfsm_g2811 : OAI221D0BWP7T port map(A1 => ml_ms_mfsm_n_17, A2 => ml_ms_mfsm_state(4), B1 => ml_ms_mfsm_state(3), B2 => ml_ms_mfsm_state(0), C => ml_ms_mfsm_n_2, ZN => ml_ms_mfsm_n_28);
  ml_ms_mfsm_g2812 : AOI22D0BWP7T port map(A1 => ml_ms_mfsm_n_18, A2 => ml_ms_mfsm_n_16, B1 => ml_ms_mfsm_n_17, B2 => ml_ms_mfsm_n_4, ZN => ml_ms_mfsm_n_27);
  ml_ms_mfsm_g2813 : MOAI22D0BWP7T port map(A1 => ml_ms_mfsm_n_20, A2 => ml_ms_mfsm_n_7, B1 => ml_ms_mfsm_n_7, B2 => ml_ms_mfsm_state(3), ZN => ml_ms_mfsm_n_26);
  ml_ms_mfsm_g2814 : IND2D1BWP7T port map(A1 => ml_ms_mfsm_n_148, B1 => ml_ms_mfsm_n_22, ZN => ml_ms_mfsm_n_25);
  ml_ms_mfsm_g2815 : ND2D1BWP7T port map(A1 => ml_ms_mfsm_n_19, A2 => ml_ms_mfsm_n_8, ZN => ml_ms_mfsm_n_24);
  ml_ms_mfsm_g2816 : OAI31D0BWP7T port map(A1 => ml_ms_count25M(10), A2 => ml_ms_count25M(9), A3 => ml_ms_mfsm_n_15, B => ml_ms_count25M(11), ZN => ml_ms_mfsm_n_23);
  ml_ms_mfsm_g2817 : INR2D1BWP7T port map(A1 => ml_ms_mfsm_n_17, B1 => ml_ms_mfsm_state(3), ZN => ml_ms_mfsm_n_21);
  ml_ms_mfsm_g2818 : NR2XD0BWP7T port map(A1 => ml_ms_mfsm_n_17, A2 => reset, ZN => ml_ms_mfsm_n_22);
  ml_ms_mfsm_g2819 : OA21D0BWP7T port map(A1 => ml_ms_mfsm_n_14, A2 => ml_ms_mfsm_state(3), B => ml_ms_mfsm_n_0, Z => ml_ms_mfsm_n_20);
  ml_ms_mfsm_g2820 : AOI222D0BWP7T port map(A1 => ml_ms_mfsm_n_9, A2 => ml_ms_mfsm_n_4, B1 => ml_ms_mfsm_n_5, B2 => ml_ms_mfsm_state(4), C1 => ml_ms_mfsm_n_3, C2 => ml_ms_mfsm_n_2, ZN => ml_ms_mfsm_n_19);
  ml_ms_mfsm_g2821 : OAI22D0BWP7T port map(A1 => ml_ms_mfsm_n_12, A2 => reset, B1 => ml_ms_mfsm_n_8, B2 => ml_ms_mfsm_state(2), ZN => ml_ms_mfsm_n_18);
  ml_ms_mfsm_g2822 : INR2XD0BWP7T port map(A1 => ml_ms_mfsm_state(0), B1 => ml_ms_mfsm_n_14, ZN => ml_ms_mfsm_n_17);
  ml_ms_mfsm_g2823 : ND2D1BWP7T port map(A1 => ml_ms_mfsm_n_14, A2 => ml_ms_mfsm_n_3, ZN => ml_ms_mfsm_n_16);
  ml_ms_mfsm_g2824 : AN4D0BWP7T port map(A1 => ml_ms_mfsm_n_6, A2 => ml_ms_count25M(8), A3 => ml_ms_count25M(6), A4 => ml_ms_count25M(7), Z => ml_ms_mfsm_n_15);
  ml_ms_mfsm_g2825 : IND2D1BWP7T port map(A1 => ml_ms_mfsm_n_10, B1 => ml_ms_count15k(3), ZN => ml_ms_mfsm_n_14);
  ml_ms_mfsm_g2826 : CKAN2D1BWP7T port map(A1 => ml_ms_mfsm_n_11, A2 => ml_ms_mfsm_n_2, Z => ml_ms_mfsm_n_13);
  ml_ms_mfsm_g2827 : ND4D0BWP7T port map(A1 => ml_ms_mfsm_n_1, A2 => ml_ms_count15k(3), A3 => ml_ms_count15k(2), A4 => ml_ms_mfsm_state(0), ZN => ml_ms_mfsm_n_12);
  ml_ms_mfsm_g2828 : AOI21D0BWP7T port map(A1 => ml_ms_count15k(0), A2 => ml_ms_count15k(1), B => ml_ms_count15k(2), ZN => ml_ms_mfsm_n_10);
  ml_ms_mfsm_g2829 : IOA21D1BWP7T port map(A1 => ml_ms_mfsm_n_148, A2 => ml_ms_mfsm_state(1), B => ml_ms_mfsm_n_0, ZN => ml_ms_mfsm_n_9);
  ml_ms_mfsm_g2830 : ND2D1BWP7T port map(A1 => ml_ms_mfsm_n_3, A2 => ml_ms_mfsm_state(0), ZN => ml_ms_mfsm_n_11);
  ml_ms_mfsm_g2831 : OR4D1BWP7T port map(A1 => ml_ms_count25M(5), A2 => ml_ms_count25M(4), A3 => ml_ms_count25M(3), A4 => ml_ms_count25M(2), Z => ml_ms_mfsm_n_6);
  ml_ms_mfsm_g2832 : ND3D0BWP7T port map(A1 => ml_ms_mfsm_state(4), A2 => ml_ms_mfsm_state(0), A3 => ml_ms_mfsm_n_2, ZN => ml_ms_mfsm_n_8);
  ml_ms_mfsm_g2833 : ND3D0BWP7T port map(A1 => ml_ms_mfsm_state(2), A2 => ml_ms_mfsm_state(0), A3 => ml_ms_mfsm_state(1), ZN => ml_ms_mfsm_n_7);
  ml_ms_mfsm_g2834 : NR2D1BWP7T port map(A1 => ml_ms_mfsm_state(1), A2 => reset, ZN => ml_ms_mfsm_n_5);
  ml_ms_mfsm_g2835 : NR2D1BWP7T port map(A1 => ml_ms_mfsm_n_1, A2 => reset, ZN => ml_ms_mfsm_n_4);
  ml_ms_mfsm_g2836 : NR2XD0BWP7T port map(A1 => ml_ms_mfsm_n_0, A2 => ml_ms_mfsm_state(3), ZN => ml_ms_mfsm_n_3);
  ml_ms_mfsm_g2837 : INVD1BWP7T port map(I => reset, ZN => ml_ms_mfsm_n_2);
  ml_ms_mfsm_state_reg_4 : DFD1BWP7T port map(CP => clk, D => ml_ms_mfsm_n_24, Q => ml_ms_mfsm_state(4), QN => ml_ms_mfsm_n_0);
  ml_ms_mfsm_state_reg_3 : DFKCND1BWP7T port map(CP => clk, CN => ml_ms_mfsm_n_2, D => ml_ms_mfsm_n_26, Q => ml_ms_mfsm_state(3), QN => ml_ms_mfsm_n_43);
  ml_ms_mfsm_state_reg_2 : DFXD1BWP7T port map(CP => clk, DA => ml_ms_mfsm_n_34, DB => ml_ms_mfsm_n_4, SA => ml_ms_mfsm_state(1), Q => ml_ms_mfsm_state(2), QN => ml_ms_mfsm_n_1);
  ml_ms_data_buffer1_Q_reg : DFQD1BWP7T port map(CP => clk, D => data_in, Q => ml_ms_Data_in_intermediate);
  ml_ms_flipflop10_Q_reg : EDFQD1BWP7T port map(CP => clk, D => ml_ms_btns(1), E => ml_ms_btnflipfloprst, Q => ml_buttons_mouse(1));
  ml_ms_flipflop1_Q_reg : EDFQD0BWP7T port map(CP => clk, D => ml_ms_mouse_x(2), E => ml_ms_xflipfloprst, Q => ml_ms_flipflop1_Q_9);
  ml_ms_flipflop1_drc_bufs : BUFFD4BWP7T port map(I => ml_ms_flipflop1_Q_9, Z => led7);
  ml_ms_data_buffer2_Q_reg : DFQD1BWP7T port map(CP => clk, D => ml_ms_Data_in_intermediate, Q => ml_ms_Data_in_buffered);
  ml_ms_tb_count_reg_3 : EDFKCNQD1BWP7T port map(CP => clk, CN => ml_ms_tb_n_1, D => ml_ms_tb_n_6, E => ml_ms_output_edgedet, Q => ml_ms_count15k(3));
  ml_ms_tb_count_reg_2 : EDFKCNQD1BWP7T port map(CP => clk, CN => ml_ms_tb_n_1, D => ml_ms_tb_n_5, E => ml_ms_output_edgedet, Q => ml_ms_count15k(2));
  ml_ms_tb_g65 : MOAI22D0BWP7T port map(A1 => ml_ms_tb_n_4, A2 => ml_ms_count15k(3), B1 => ml_ms_tb_n_4, B2 => ml_ms_count15k(3), ZN => ml_ms_tb_n_6);
  ml_ms_tb_count_reg_1 : EDFKCNQD1BWP7T port map(CP => clk, CN => ml_ms_tb_n_1, D => ml_ms_tb_n_3, E => ml_ms_output_edgedet, Q => ml_ms_count15k(1));
  ml_ms_tb_g67 : MOAI22D0BWP7T port map(A1 => ml_ms_tb_n_2, A2 => ml_ms_count15k(2), B1 => ml_ms_tb_n_2, B2 => ml_ms_count15k(2), ZN => ml_ms_tb_n_5);
  ml_ms_tb_count_reg_0 : DFKCNQD1BWP7T port map(CP => clk, CN => ml_ms_tb_n_0, D => ml_ms_tb_n_1, Q => ml_ms_count15k(0));
  ml_ms_tb_g69 : IND2D1BWP7T port map(A1 => ml_ms_tb_n_2, B1 => ml_ms_count15k(2), ZN => ml_ms_tb_n_4);
  ml_ms_tb_g70 : CKXOR2D0BWP7T port map(A1 => ml_ms_count15k(1), A2 => ml_ms_count15k(0), Z => ml_ms_tb_n_3);
  ml_ms_tb_g72 : ND2D1BWP7T port map(A1 => ml_ms_count15k(1), A2 => ml_ms_count15k(0), ZN => ml_ms_tb_n_2);
  ml_ms_tb_g73 : INVD1BWP7T port map(I => ml_ms_cntReset15K, ZN => ml_ms_tb_n_1);
  ml_ms_tb_g2 : CKXOR2D1BWP7T port map(A1 => ml_ms_output_edgedet, A2 => ml_ms_count15k(0), Z => ml_ms_tb_n_0);
  ml_ms_flipflop11_Q_reg : EDFQD1BWP7T port map(CP => clk, D => ml_ms_btns(0), E => ml_ms_btnflipfloprst, Q => ml_ms_n_82);
  ml_ms_flipflop2_Q_reg : EDFQD1BWP7T port map(CP => clk, D => ml_ms_mouse_x(1), E => ml_ms_xflipfloprst, Q => ml_mouseX(1));
  ml_ms_sr11_g27 : INVD1BWP7T port map(I => reset, ZN => ml_ms_sr11_n_0);
  ml_ms_sr11_data_out_reg_3 : EDFKCNQD1BWP7T port map(CP => clk, CN => ml_ms_sr11_n_0, D => ml_ms_sr11_data_out_2_81, E => ml_ms_output_edgedet, Q => ml_ms_sr11_data_out_3_82);
  ml_ms_sr11_data_out_reg_1 : EDFKCNQD1BWP7T port map(CP => clk, CN => ml_ms_sr11_n_0, D => ml_ms_sr11_data_out_0_79, E => ml_ms_output_edgedet, Q => ml_ms_sr11_data_out_1_80);
  ml_ms_sr11_data_out_reg_0 : EDFKCNQD1BWP7T port map(CP => clk, CN => ml_ms_sr11_n_0, D => ml_ms_Data_in_buffered, E => ml_ms_output_edgedet, Q => ml_ms_sr11_data_out_0_79);
  ml_ms_sr11_data_out_reg_9 : EDFKCNQD1BWP7T port map(CP => clk, CN => ml_ms_sr11_n_0, D => ml_ms_data_sr_11bit(8), E => ml_ms_output_edgedet, Q => ml_ms_data_sr_11bit(9));
  ml_ms_sr11_data_out_reg_4 : EDFKCNQD1BWP7T port map(CP => clk, CN => ml_ms_sr11_n_0, D => ml_ms_sr11_data_out_3_82, E => ml_ms_output_edgedet, Q => ml_ms_data_sr_11bit(4));
  ml_ms_sr11_data_out_reg_2 : EDFKCNQD1BWP7T port map(CP => clk, CN => ml_ms_sr11_n_0, D => ml_ms_sr11_data_out_1_80, E => ml_ms_output_edgedet, Q => ml_ms_sr11_data_out_2_81);
  ml_ms_sr11_data_out_reg_6 : EDFKCNQD1BWP7T port map(CP => clk, CN => ml_ms_sr11_n_0, D => ml_ms_data_sr_11bit(5), E => ml_ms_output_edgedet, Q => ml_ms_data_sr_11bit(6));
  ml_ms_sr11_data_out_reg_5 : EDFKCNQD1BWP7T port map(CP => clk, CN => ml_ms_sr11_n_0, D => ml_ms_data_sr_11bit(4), E => ml_ms_output_edgedet, Q => ml_ms_data_sr_11bit(5));
  ml_ms_sr11_data_out_reg_7 : EDFKCNQD1BWP7T port map(CP => clk, CN => ml_ms_sr11_n_0, D => ml_ms_data_sr_11bit(6), E => ml_ms_output_edgedet, Q => ml_ms_data_sr_11bit(7));
  ml_ms_sr11_data_out_reg_8 : EDFKCNQD1BWP7T port map(CP => clk, CN => ml_ms_sr11_n_0, D => ml_ms_data_sr_11bit(7), E => ml_ms_output_edgedet, Q => ml_ms_data_sr_11bit(8));
  ml_ms_flipflop3_Q_reg : EDFQD1BWP7T port map(CP => clk, D => ml_ms_mouse_x(0), E => ml_ms_xflipfloprst, Q => ml_ms_n_78);
  ml_ms_flipflop4_Q_reg : EDFQD1BWP7T port map(CP => clk, D => ml_ms_mouse_y(0), E => ml_ms_yflipfloprst, Q => ml_ms_flipflop4_Q_9);
  ml_ms_flipflop4_drc_bufs : BUFFD4BWP7T port map(I => ml_ms_flipflop4_Q_9, Z => led3);
  ml_il_y1_tempy_reg_2 : DFQD1BWP7T port map(CP => clk, D => ml_il_y1_n_28, Q => sig_logic_y(2));
  ml_il_y1_g635 : OR2D1BWP7T port map(A1 => ml_il_y1_locy(2), A2 => reset, Z => ml_il_y1_n_28);
  ml_il_y1_tempy_reg_1 : DFKCNQD1BWP7T port map(CP => clk, CN => ml_il_y1_n_0, D => ml_il_y1_locy(1), Q => sig_logic_y(1));
  ml_il_y1_tempy_reg_0 : DFKSND1BWP7T port map(CP => clk, D => ml_il_y1_locy(0), SN => ml_il_y1_n_0, Q => sig_logic_y(0), QN => UNCONNECTED);
  ml_il_y1_g638 : OR3D1BWP7T port map(A1 => ml_il_y1_n_25, A2 => ml_il_y1_n_32, A3 => ml_il_y1_n_27, Z => ml_il_y1_locy(2));
  ml_il_y1_g639 : OR4D1BWP7T port map(A1 => ml_il_y1_n_12, A2 => ml_il_y1_n_14, A3 => ml_il_y1_n_25, A4 => ml_il_y1_n_32, Z => ml_il_y1_locy(0));
  ml_il_y1_g640 : AO22D0BWP7T port map(A1 => ml_il_y1_n_33, A2 => ml_il_y1_n_22, B1 => ml_il_y1_n_23, B2 => ml_il_y1_n_31, Z => ml_il_y1_n_27);
  ml_il_y1_g641 : AO22D0BWP7T port map(A1 => ml_il_y1_n_33, A2 => ml_il_y1_n_41, B1 => ml_il_y1_n_20, B2 => ml_il_y1_n_31, Z => ml_il_y1_locy(1));
  ml_il_y1_g642 : AN2D1BWP7T port map(A1 => ml_il_y1_n_26, A2 => ml_buttons_mouse(1), Z => ml_il_y1_n_33);
  ml_il_y1_g643 : INR2D1BWP7T port map(A1 => ml_buttons_mouse(1), B1 => ml_il_y1_n_26, ZN => ml_il_y1_n_32);
  ml_il_y1_g644 : OAI211D1BWP7T port map(A1 => ml_il_y1_input_register(1), A2 => ml_il_y1_n_18, B => ml_il_y1_n_24, C => ml_il_y1_input_register(3), ZN => ml_il_y1_n_26);
  ml_il_y1_g645 : AOI21D0BWP7T port map(A1 => ml_il_y1_n_40, A2 => ml_il_y1_n_29, B => ml_buttons_mouse(1), ZN => ml_il_y1_n_31);
  ml_il_y1_g646 : INR3D0BWP7T port map(A1 => ml_il_y1_n_40, B1 => ml_il_y1_input_register(3), B2 => ml_buttons_mouse(1), ZN => ml_il_y1_n_25);
  ml_il_y1_g647 : AO21D0BWP7T port map(A1 => ml_il_y1_n_18, A2 => ml_il_y1_input_register(1), B => ml_il_y1_input_register(2), Z => ml_il_y1_n_24);
  ml_il_y1_g648 : MOAI22D0BWP7T port map(A1 => ml_il_y1_n_36, A2 => ml_il_y1_input_register(2), B1 => ml_il_y1_n_36, B2 => ml_il_y1_input_register(2), ZN => ml_il_y1_n_23);
  ml_il_y1_g649 : MOAI22D0BWP7T port map(A1 => ml_il_y1_n_30, A2 => ml_il_y1_n_39, B1 => ml_il_y1_n_30, B2 => ml_il_y1_n_39, ZN => ml_il_y1_n_22);
  ml_il_y1_g651 : MOAI22D0BWP7T port map(A1 => ml_il_y1_n_17, A2 => ml_il_y1_n_12, B1 => ml_il_y1_n_17, B2 => ml_il_y1_n_12, ZN => ml_il_y1_n_20);
  ml_il_y1_g653 : AOI21D0BWP7T port map(A1 => ml_il_y1_n_8, A2 => ml_il_y1_n_7, B => ml_il_y1_n_9, ZN => ml_il_y1_n_18);
  ml_il_y1_g654 : OAI21D0BWP7T port map(A1 => ml_il_y1_n_13, A2 => ml_il_y1_n_7, B => ml_il_y1_n_10, ZN => ml_il_y1_n_30);
  ml_il_y1_g655 : AO21D0BWP7T port map(A1 => ml_il_y1_n_8, A2 => ml_il_y1_n_11, B => ml_il_y1_n_9, Z => ml_il_y1_n_36);
  ml_il_y1_g657 : IND2D1BWP7T port map(A1 => ml_il_y1_n_13, B1 => ml_il_y1_n_10, ZN => ml_il_y1_n_17);
  ml_il_y1_g659 : INVD0BWP7T port map(I => ml_il_y1_n_11, ZN => ml_il_y1_n_12);
  ml_il_y1_g660 : INR2D1BWP7T port map(A1 => ml_il_y1_input_register(0), B1 => led3, ZN => ml_il_y1_n_14);
  ml_il_y1_g661 : NR2XD0BWP7T port map(A1 => led2, A2 => ml_il_y1_input_register(1), ZN => ml_il_y1_n_13);
  ml_il_y1_g662 : IND2D1BWP7T port map(A1 => ml_il_y1_input_register(0), B1 => led3, ZN => ml_il_y1_n_11);
  ml_il_y1_g663 : ND2D1BWP7T port map(A1 => led2, A2 => ml_il_y1_input_register(1), ZN => ml_il_y1_n_10);
  ml_il_y1_g664 : INR2D1BWP7T port map(A1 => ml_il_y1_input_register(1), B1 => led2, ZN => ml_il_y1_n_9);
  ml_il_y1_g665 : IND2D1BWP7T port map(A1 => ml_il_y1_input_register(1), B1 => led2, ZN => ml_il_y1_n_8);
  ml_il_y1_g666 : ND2D1BWP7T port map(A1 => led3, A2 => ml_il_y1_input_register(0), ZN => ml_il_y1_n_7);
  ml_il_y1_g668 : INVD0BWP7T port map(I => reset, ZN => ml_il_y1_n_0);
  ml_il_y1_tempy_reg_3 : DFKCNQD1BWP7T port map(CP => clk, CN => ml_il_y1_n_0, D => ml_il_y1_n_5, Q => sig_logic_y(3));
  ml_il_y1_g333 : AO221D0BWP7T port map(A1 => ml_il_y1_n_4, A2 => ml_il_y1_n_31, B1 => ml_il_y1_n_33, B2 => ml_il_y1_n_3, C => ml_il_y1_n_32, Z => ml_il_y1_n_5);
  ml_il_y1_input_register_reg_0 : DFXQD1BWP7T port map(CP => clk, DA => ml_il_y1_locy(0), DB => sig_logic_y(0), SA => ml_handshake_mouse_out, Q => ml_il_y1_input_register(0));
  ml_il_y1_input_register_reg_1 : DFXQD1BWP7T port map(CP => clk, DA => ml_il_y1_locy(1), DB => sig_logic_y(1), SA => ml_handshake_mouse_out, Q => ml_il_y1_input_register(1));
  ml_il_y1_g337 : MOAI22D0BWP7T port map(A1 => ml_il_y1_n_2, A2 => ml_il_y1_input_register(3), B1 => ml_il_y1_n_2, B2 => ml_il_y1_input_register(3), ZN => ml_il_y1_n_4);
  ml_il_y1_g338 : MOAI22D0BWP7T port map(A1 => ml_il_y1_n_1, A2 => ml_il_y1_n_29, B1 => ml_il_y1_n_1, B2 => ml_il_y1_n_29, ZN => ml_il_y1_n_3);
  ml_il_y1_g339 : IND2D1BWP7T port map(A1 => ml_il_y1_n_36, B1 => ml_il_y1_n_39, ZN => ml_il_y1_n_2);
  ml_il_y1_g340 : AN2D0BWP7T port map(A1 => ml_il_y1_n_30, A2 => ml_il_y1_input_register(2), Z => ml_il_y1_n_1);
  ml_il_y1_g2 : ND2D1BWP7T port map(A1 => ml_il_y1_n_9, A2 => ml_il_y1_input_register(2), ZN => ml_il_y1_n_40);
  ml_il_y1_g670 : CKXOR2D1BWP7T port map(A1 => ml_il_y1_n_17, A2 => ml_il_y1_n_7, Z => ml_il_y1_n_41);
  ml_il_y1_input_register_reg_3 : DFXD1BWP7T port map(CP => clk, DA => ml_il_y1_n_5, DB => sig_logic_y(3), SA => ml_handshake_mouse_out, Q => ml_il_y1_input_register(3), QN => ml_il_y1_n_29);
  ml_il_y1_input_register_reg_2 : DFXD1BWP7T port map(CP => clk, DA => ml_il_y1_locy(2), DB => sig_logic_y(2), SA => ml_handshake_mouse_out, Q => ml_il_y1_input_register(2), QN => ml_il_y1_n_39);
  ml_ms_flipflop5_Q_reg : EDFQD1BWP7T port map(CP => clk, D => ml_ms_mouse_y(1), E => ml_ms_yflipfloprst, Q => ml_ms_flipflop5_Q_9);
  ml_ms_flipflop5_drc_bufs : BUFFD4BWP7T port map(I => ml_ms_flipflop5_Q_9, Z => led2);
  ml_ms_flipflop6_Q_reg : EDFQD0BWP7T port map(CP => clk, D => ml_ms_mouse_y(2), E => ml_ms_yflipfloprst, Q => ml_ms_flipflop6_Q_9);
  ml_ms_flipflop6_drc_bufs : BUFFD4BWP7T port map(I => ml_ms_flipflop6_Q_9, Z => led1);
  ml_ms_flipflop7_Q_reg : EDFQD1BWP7T port map(CP => clk, D => ml_ms_btns(4), E => ml_ms_btnflipfloprst, Q => ml_buttons_mouse(4));
  ml_ms_flipflop8_Q_reg : DFXQD1BWP7T port map(CP => clk, DA => ml_ms_btns(3), DB => sig_middelsteknop, SA => ml_ms_btnflipfloprst, Q => sig_middelsteknop);
  ml_ms_clk_buffer1_Q_reg : DFQD1BWP7T port map(CP => clk, D => clk15k_in, Q => ml_ms_Clk15k_intermediate);
  ml_ms_mx_g23 : ND2D4BWP7T port map(A1 => ml_ms_mx_n_0, A2 => ml_ms_mx_n_1, ZN => data_switch);
  ml_ms_mx_g24 : ND2D1BWP7T port map(A1 => ml_ms_mux_select, A2 => ml_ms_muxReg, ZN => ml_ms_mx_n_1);
  ml_ms_mx_g25 : IND2D1BWP7T port map(A1 => ml_ms_mux_select, B1 => ml_ms_muxFSM, ZN => ml_ms_mx_n_0);
  ml_ms_flipflop9_Q_reg : EDFQD1BWP7T port map(CP => clk, D => ml_ms_btns(2), E => ml_ms_btnflipfloprst, Q => sig_draw);
  ml_ms_cnt_g71 : CKND1BWP7T port map(I => ml_ms_cntReset25M, ZN => ml_ms_cnt_n_23);
  ml_ms_cnt_count_reg_12 : DFKCNQD1BWP7T port map(CP => clk, CN => ml_ms_cnt_n_23, D => ml_ms_cnt_n_22, Q => ml_ms_count25M(12));
  ml_ms_cnt_count_reg_11 : DFKCNQD1BWP7T port map(CP => clk, CN => ml_ms_cnt_n_23, D => ml_ms_cnt_n_21, Q => ml_ms_count25M(11));
  ml_ms_cnt_g225 : MOAI22D0BWP7T port map(A1 => ml_ms_cnt_n_20, A2 => ml_ms_count25M(12), B1 => ml_ms_cnt_n_20, B2 => ml_ms_count25M(12), ZN => ml_ms_cnt_n_22);
  ml_ms_cnt_count_reg_10 : DFKCNQD1BWP7T port map(CP => clk, CN => ml_ms_cnt_n_23, D => ml_ms_cnt_n_19, Q => ml_ms_count25M(10));
  ml_ms_cnt_g227 : MOAI22D0BWP7T port map(A1 => ml_ms_cnt_n_18, A2 => ml_ms_count25M(11), B1 => ml_ms_cnt_n_18, B2 => ml_ms_count25M(11), ZN => ml_ms_cnt_n_21);
  ml_ms_cnt_g228 : IND2D1BWP7T port map(A1 => ml_ms_cnt_n_18, B1 => ml_ms_count25M(11), ZN => ml_ms_cnt_n_20);
  ml_ms_cnt_count_reg_9 : DFKCNQD1BWP7T port map(CP => clk, CN => ml_ms_cnt_n_23, D => ml_ms_cnt_n_17, Q => ml_ms_count25M(9));
  ml_ms_cnt_g230 : MOAI22D0BWP7T port map(A1 => ml_ms_cnt_n_16, A2 => ml_ms_count25M(10), B1 => ml_ms_cnt_n_16, B2 => ml_ms_count25M(10), ZN => ml_ms_cnt_n_19);
  ml_ms_cnt_g231 : IND2D1BWP7T port map(A1 => ml_ms_cnt_n_16, B1 => ml_ms_count25M(10), ZN => ml_ms_cnt_n_18);
  ml_ms_cnt_count_reg_8 : DFKCNQD1BWP7T port map(CP => clk, CN => ml_ms_cnt_n_23, D => ml_ms_cnt_n_15, Q => ml_ms_count25M(8));
  ml_ms_cnt_g233 : MOAI22D0BWP7T port map(A1 => ml_ms_cnt_n_14, A2 => ml_ms_count25M(9), B1 => ml_ms_cnt_n_14, B2 => ml_ms_count25M(9), ZN => ml_ms_cnt_n_17);
  ml_ms_cnt_g234 : IND2D1BWP7T port map(A1 => ml_ms_cnt_n_14, B1 => ml_ms_count25M(9), ZN => ml_ms_cnt_n_16);
  ml_ms_cnt_count_reg_7 : DFKCNQD1BWP7T port map(CP => clk, CN => ml_ms_cnt_n_23, D => ml_ms_cnt_n_13, Q => ml_ms_count25M(7));
  ml_ms_cnt_g236 : MOAI22D0BWP7T port map(A1 => ml_ms_cnt_n_12, A2 => ml_ms_count25M(8), B1 => ml_ms_cnt_n_12, B2 => ml_ms_count25M(8), ZN => ml_ms_cnt_n_15);
  ml_ms_cnt_g237 : IND2D1BWP7T port map(A1 => ml_ms_cnt_n_12, B1 => ml_ms_count25M(8), ZN => ml_ms_cnt_n_14);
  ml_ms_cnt_count_reg_6 : DFKCNQD1BWP7T port map(CP => clk, CN => ml_ms_cnt_n_11, D => ml_ms_cnt_n_23, Q => ml_ms_count25M(6));
  ml_ms_cnt_g239 : MOAI22D0BWP7T port map(A1 => ml_ms_cnt_n_10, A2 => ml_ms_count25M(7), B1 => ml_ms_cnt_n_10, B2 => ml_ms_count25M(7), ZN => ml_ms_cnt_n_13);
  ml_ms_cnt_g240 : IND2D1BWP7T port map(A1 => ml_ms_cnt_n_10, B1 => ml_ms_count25M(7), ZN => ml_ms_cnt_n_12);
  ml_ms_cnt_count_reg_5 : DFKCNQD1BWP7T port map(CP => clk, CN => ml_ms_cnt_n_9, D => ml_ms_cnt_n_23, Q => ml_ms_count25M(5));
  ml_ms_cnt_g242 : MOAI22D0BWP7T port map(A1 => ml_ms_cnt_n_8, A2 => ml_ms_count25M(6), B1 => ml_ms_cnt_n_8, B2 => ml_ms_count25M(6), ZN => ml_ms_cnt_n_11);
  ml_ms_cnt_g243 : IND2D1BWP7T port map(A1 => ml_ms_cnt_n_8, B1 => ml_ms_count25M(6), ZN => ml_ms_cnt_n_10);
  ml_ms_cnt_count_reg_4 : DFKCNQD1BWP7T port map(CP => clk, CN => ml_ms_cnt_n_7, D => ml_ms_cnt_n_23, Q => ml_ms_count25M(4));
  ml_ms_cnt_g245 : MOAI22D0BWP7T port map(A1 => ml_ms_cnt_n_6, A2 => ml_ms_count25M(5), B1 => ml_ms_cnt_n_6, B2 => ml_ms_count25M(5), ZN => ml_ms_cnt_n_9);
  ml_ms_cnt_g246 : IND2D1BWP7T port map(A1 => ml_ms_cnt_n_6, B1 => ml_ms_count25M(5), ZN => ml_ms_cnt_n_8);
  ml_ms_cnt_count_reg_3 : DFKCNQD1BWP7T port map(CP => clk, CN => ml_ms_cnt_n_5, D => ml_ms_cnt_n_23, Q => ml_ms_count25M(3));
  ml_ms_cnt_g248 : MOAI22D0BWP7T port map(A1 => ml_ms_cnt_n_4, A2 => ml_ms_count25M(4), B1 => ml_ms_cnt_n_4, B2 => ml_ms_count25M(4), ZN => ml_ms_cnt_n_7);
  ml_ms_cnt_g249 : IND2D1BWP7T port map(A1 => ml_ms_cnt_n_4, B1 => ml_ms_count25M(4), ZN => ml_ms_cnt_n_6);
  ml_ms_cnt_count_reg_2 : DFKCNQD1BWP7T port map(CP => clk, CN => ml_ms_cnt_n_3, D => ml_ms_cnt_n_23, Q => ml_ms_count25M(2));
  ml_ms_cnt_g251 : MOAI22D0BWP7T port map(A1 => ml_ms_cnt_n_2, A2 => ml_ms_count25M(3), B1 => ml_ms_cnt_n_2, B2 => ml_ms_count25M(3), ZN => ml_ms_cnt_n_5);
  ml_ms_cnt_g252 : IND2D1BWP7T port map(A1 => ml_ms_cnt_n_2, B1 => ml_ms_count25M(3), ZN => ml_ms_cnt_n_4);
  ml_ms_cnt_count_reg_1 : EDFKCND1BWP7T port map(CP => clk, CN => ml_ms_cnt_n_23, D => ml_ms_cnt_count(1), E => ml_ms_cnt_count(0), Q => UNCONNECTED0, QN => ml_ms_cnt_count(1));
  ml_ms_cnt_g254 : MOAI22D0BWP7T port map(A1 => ml_ms_cnt_n_1, A2 => ml_ms_count25M(2), B1 => ml_ms_cnt_n_1, B2 => ml_ms_count25M(2), ZN => ml_ms_cnt_n_3);
  ml_ms_cnt_g255 : IND2D1BWP7T port map(A1 => ml_ms_cnt_n_1, B1 => ml_ms_count25M(2), ZN => ml_ms_cnt_n_2);
  ml_ms_cnt_g257 : IND2D1BWP7T port map(A1 => ml_ms_cnt_count(1), B1 => ml_ms_cnt_count(0), ZN => ml_ms_cnt_n_1);
  ml_ms_cnt_count_reg_0 : DFKCND1BWP7T port map(CP => clk, CN => ml_ms_cnt_n_0, D => ml_ms_cnt_n_23, Q => ml_ms_cnt_count(0), QN => ml_ms_cnt_n_0);
  ml_ms_clk_buffer2_Q_reg : DFQD1BWP7T port map(CP => clk, D => ml_ms_Clk15k_intermediate, Q => ml_ms_Clk15k_buffered);
  ml_il_color1_g570 : AO21D0BWP7T port map(A1 => sig_output_color(1), A2 => ml_il_color1_n_16, B => ml_il_color1_n_22, Z => sig_output_color(0));
  ml_il_color1_g571 : HA1D0BWP7T port map(A => ml_il_color1_state(2), B => ml_il_color1_state(1), CO => ml_il_color1_n_22, S => sig_output_color(1));
  ml_il_color1_g572 : OAI21D0BWP7T port map(A1 => ml_il_color1_n_17, A2 => ml_il_color1_state(1), B => ml_il_color1_n_23, ZN => sig_output_color(2));
  ml_il_color1_g573 : ND2D1BWP7T port map(A1 => ml_il_color1_state(0), A2 => ml_il_color1_state(2), ZN => ml_il_color1_n_23);
  ml_il_color1_g574 : NR2D0BWP7T port map(A1 => ml_il_color1_state(0), A2 => ml_il_color1_state(2), ZN => ml_il_color1_n_17);
  ml_il_color1_state_reg_1 : DFKSND1BWP7T port map(CP => clk, D => reset, SN => ml_il_color1_n_15, Q => ml_il_color1_state(1), QN => ml_il_color1_n_0);
  ml_il_color1_state_reg_2 : DFKCNQD1BWP7T port map(CP => clk, CN => ml_il_color1_n_9, D => ml_il_color1_n_14, Q => ml_il_color1_state(2));
  ml_il_color1_g805 : INR4D0BWP7T port map(A1 => ml_il_color1_n_9, B1 => ml_il_color1_n_22, B2 => ml_il_color1_n_7, B3 => ml_il_color1_n_12, ZN => ml_il_color1_n_15);
  ml_il_color1_state_hs_reg_1 : DFKCNQD1BWP7T port map(CP => clk, CN => ml_il_color1_n_1, D => ml_il_color1_n_10, Q => ml_il_color1_state_hs(1));
  ml_il_color1_g808 : OAI211D1BWP7T port map(A1 => ml_il_color1_n_0, A2 => ml_il_color1_n_7, B => ml_il_color1_n_11, C => ml_il_color1_n_1, ZN => ml_il_color1_n_14);
  ml_il_color1_g809 : AO21D0BWP7T port map(A1 => ml_il_color1_n_8, A2 => ml_il_color1_n_1, B => ml_il_color1_n_5, Z => ml_il_color1_n_13);
  ml_il_color1_state_hs_reg_0 : DFKCNQD1BWP7T port map(CP => clk, CN => ml_il_color1_n_6, D => ml_handshake_mouse_out, Q => ml_il_color1_state_hs(0));
  ml_il_color1_g811 : AN3D0BWP7T port map(A1 => ml_il_color1_n_5, A2 => ml_il_color1_n_2, A3 => ml_il_color1_n_0, Z => ml_il_color1_n_12);
  ml_il_color1_g812 : OAI21D0BWP7T port map(A1 => ml_il_color1_n_3, A2 => ml_il_color1_n_4, B => ml_il_color1_state(2), ZN => ml_il_color1_n_11);
  ml_il_color1_g813 : IAO21D0BWP7T port map(A1 => ml_handshake_mouse_out, A2 => ml_il_color1_state_hs(0), B => ml_il_color1_n_6, ZN => ml_il_color1_n_10);
  ml_il_color1_g814 : OAI32D1BWP7T port map(A1 => ml_il_color1_state(0), A2 => ml_il_color1_n_3, A3 => sig_output_color(1), B1 => ml_il_color1_n_23, B2 => ml_il_color1_n_2, ZN => ml_il_color1_n_8);
  ml_il_color1_g815 : IND4D0BWP7T port map(A1 => ml_il_color1_state(2), B1 => ml_il_color1_n_1, B2 => ml_il_color1_state(1), B3 => ml_il_color1_n_3, ZN => ml_il_color1_n_9);
  ml_il_color1_g816 : NR2D1BWP7T port map(A1 => ml_il_color1_n_23, A2 => ml_il_color1_n_3, ZN => ml_il_color1_n_7);
  ml_il_color1_g817 : NR3D0BWP7T port map(A1 => ml_il_color1_state_hs(0), A2 => ml_il_color1_state_hs(1), A3 => reset, ZN => ml_il_color1_n_6);
  ml_il_color1_g818 : INR3D0BWP7T port map(A1 => ml_il_color1_state(0), B1 => reset, B2 => ml_il_color1_state(2), ZN => ml_il_color1_n_5);
  ml_il_color1_g819 : AN2D0BWP7T port map(A1 => ml_il_color1_n_0, A2 => ml_il_color1_state(0), Z => ml_il_color1_n_4);
  ml_il_color1_g820 : INVD0BWP7T port map(I => ml_il_color1_n_3, ZN => ml_il_color1_n_2);
  ml_il_color1_g821 : ND2D1BWP7T port map(A1 => ml_buttons_mouse(4), A2 => ml_il_color1_state_hs(0), ZN => ml_il_color1_n_3);
  ml_il_color1_g826 : INVD1BWP7T port map(I => reset, ZN => ml_il_color1_n_1);
  ml_il_color1_state_reg_0 : DFD1BWP7T port map(CP => clk, D => ml_il_color1_n_13, Q => ml_il_color1_state(0), QN => ml_il_color1_n_16);
  ml_il_x1_tempx_reg_0 : DFQD1BWP7T port map(CP => clk, D => ml_il_x1_n_25, Q => sig_logic_x(0));
  ml_il_x1_tempx_reg_1 : DFQD1BWP7T port map(CP => clk, D => ml_il_x1_n_24, Q => sig_logic_x(1));
  ml_il_x1_tempx_reg_3 : DFQD1BWP7T port map(CP => clk, D => ml_il_x1_n_23, Q => sig_logic_x(3));
  ml_il_x1_g634 : AO211D0BWP7T port map(A1 => ml_il_x1_n_18, A2 => led6, B => ml_il_x1_n_22, C => reset, Z => ml_il_x1_n_25);
  ml_il_x1_g635 : AO221D0BWP7T port map(A1 => ml_il_x1_n_28, A2 => ml_il_x1_n_14, B1 => ml_il_x1_n_29, B2 => ml_il_x1_n_15, C => ml_il_x1_n_21, Z => ml_il_x1_n_24);
  ml_il_x1_g636 : AO221D0BWP7T port map(A1 => ml_il_x1_n_20, A2 => ml_il_x1_input_register(3), B1 => ml_il_x1_n_29, B2 => ml_il_x1_n_17, C => ml_il_x1_n_21, Z => ml_il_x1_n_23);
  ml_il_x1_g637 : MAOI22D0BWP7T port map(A1 => ml_il_x1_n_7, A2 => ml_il_x1_n_9, B1 => ml_il_x1_n_28, B2 => ml_il_x1_n_29, ZN => ml_il_x1_n_22);
  ml_il_x1_g638 : NR3D0BWP7T port map(A1 => ml_il_x1_n_19, A2 => led6, A3 => reset, ZN => ml_il_x1_n_21);
  ml_il_x1_g639 : OA21D0BWP7T port map(A1 => ml_il_x1_n_26, A2 => ml_il_x1_input_register(2), B => ml_il_x1_n_28, Z => ml_il_x1_n_20);
  ml_il_x1_g640 : INR3D0BWP7T port map(A1 => ml_il_x1_n_19, B1 => reset, B2 => led6, ZN => ml_il_x1_n_29);
  ml_il_x1_g641 : INR3D0BWP7T port map(A1 => led6, B1 => reset, B2 => ml_il_x1_n_18, ZN => ml_il_x1_n_28);
  ml_il_x1_g642 : OAI21D0BWP7T port map(A1 => ml_il_x1_n_16, A2 => ml_il_x1_input_register(2), B => ml_il_x1_input_register(3), ZN => ml_il_x1_n_19);
  ml_il_x1_g643 : NR4D0BWP7T port map(A1 => ml_il_x1_n_12, A2 => ml_il_x1_n_11, A3 => ml_il_x1_input_register(3), A4 => ml_il_x1_input_register(2), ZN => ml_il_x1_n_18);
  ml_il_x1_g644 : AO21D0BWP7T port map(A1 => ml_il_x1_n_27, A2 => ml_il_x1_input_register(2), B => ml_il_x1_input_register(3), Z => ml_il_x1_n_17);
  ml_il_x1_g645 : OA31D1BWP7T port map(A1 => ml_il_x1_input_register(0), A2 => led9, A3 => ml_il_x1_n_10, B => ml_il_x1_n_6, Z => ml_il_x1_n_16);
  ml_il_x1_g646 : MOAI22D0BWP7T port map(A1 => ml_il_x1_n_13, A2 => ml_il_x1_n_5, B1 => ml_il_x1_n_13, B2 => ml_il_x1_n_5, ZN => ml_il_x1_n_15);
  ml_il_x1_g647 : MOAI22D0BWP7T port map(A1 => ml_il_x1_n_13, A2 => ml_il_x1_n_9, B1 => ml_il_x1_n_13, B2 => ml_il_x1_n_9, ZN => ml_il_x1_n_14);
  ml_il_x1_g648 : AO21D0BWP7T port map(A1 => ml_il_x1_n_6, A2 => ml_il_x1_n_4, B => ml_il_x1_n_10, Z => ml_il_x1_n_27);
  ml_il_x1_g649 : AO21D0BWP7T port map(A1 => ml_il_x1_n_8, A2 => ml_il_x1_n_9, B => ml_il_x1_n_11, Z => ml_il_x1_n_26);
  ml_il_x1_g650 : INR2D1BWP7T port map(A1 => ml_il_x1_n_6, B1 => ml_il_x1_n_10, ZN => ml_il_x1_n_13);
  ml_il_x1_g651 : INR2D1BWP7T port map(A1 => ml_il_x1_n_8, B1 => ml_il_x1_n_7, ZN => ml_il_x1_n_12);
  ml_il_x1_g652 : INR2D1BWP7T port map(A1 => ml_il_x1_input_register(1), B1 => ml_mouseX(1), ZN => ml_il_x1_n_11);
  ml_il_x1_g653 : AN2D1BWP7T port map(A1 => ml_il_x1_input_register(1), A2 => ml_mouseX(1), Z => ml_il_x1_n_10);
  ml_il_x1_g654 : IND2D1BWP7T port map(A1 => ml_il_x1_input_register(0), B1 => led9, ZN => ml_il_x1_n_9);
  ml_il_x1_input_register_reg_2 : DFQD1BWP7T port map(CP => clk, D => sig_logic_x(2), Q => ml_il_x1_input_register(2));
  ml_il_x1_g656 : INVD1BWP7T port map(I => ml_il_x1_n_5, ZN => ml_il_x1_n_4);
  ml_il_x1_g657 : IND2D1BWP7T port map(A1 => ml_il_x1_input_register(1), B1 => ml_mouseX(1), ZN => ml_il_x1_n_8);
  ml_il_x1_g658 : IND2D1BWP7T port map(A1 => led9, B1 => ml_il_x1_input_register(0), ZN => ml_il_x1_n_7);
  ml_il_x1_g659 : OR2D1BWP7T port map(A1 => ml_il_x1_input_register(1), A2 => ml_mouseX(1), Z => ml_il_x1_n_6);
  ml_il_x1_g660 : ND2D1BWP7T port map(A1 => led9, A2 => ml_il_x1_input_register(0), ZN => ml_il_x1_n_5);
  ml_il_x1_tempx_reg_2 : DFXQD1BWP7T port map(CP => clk, DA => ml_il_x1_n_3, DB => ml_il_x1_n_2, SA => ml_il_x1_input_register(2), Q => sig_logic_x(2));
  ml_il_x1_g277 : MOAI22D0BWP7T port map(A1 => ml_il_x1_n_0, A2 => ml_il_x1_n_27, B1 => ml_il_x1_n_28, B2 => ml_il_x1_n_26, ZN => ml_il_x1_n_3);
  ml_il_x1_g278 : MOAI22D0BWP7T port map(A1 => ml_il_x1_n_1, A2 => ml_il_x1_n_26, B1 => ml_il_x1_n_29, B2 => ml_il_x1_n_27, ZN => ml_il_x1_n_2);
  ml_il_x1_input_register_reg_0 : DFQD1BWP7T port map(CP => clk, D => sig_logic_x(0), Q => ml_il_x1_input_register(0));
  ml_il_x1_input_register_reg_1 : DFQD1BWP7T port map(CP => clk, D => sig_logic_x(1), Q => ml_il_x1_input_register(1));
  ml_il_x1_input_register_reg_3 : DFQD1BWP7T port map(CP => clk, D => sig_logic_x(3), Q => ml_il_x1_input_register(3));
  ml_il_x1_g282 : INVD0BWP7T port map(I => ml_il_x1_n_28, ZN => ml_il_x1_n_1);
  ml_il_x1_g283 : INVD0BWP7T port map(I => ml_il_x1_n_29, ZN => ml_il_x1_n_0);
  gl_vgd_g1606 : OR2D4BWP7T port map(A1 => gl_vgd_n_81, A2 => gl_vgd_horizontal(8), Z => H);
  gl_vgd_g1607 : ND2D1BWP7T port map(A1 => gl_vgd_n_80, A2 => gl_vgd_horizontal(9), ZN => gl_vgd_n_81);
  gl_vgd_g1608 : AN2D4BWP7T port map(A1 => gl_sig_red, A2 => gl_vgd_n_79, Z => R);
  gl_vgd_g1609 : AN2D4BWP7T port map(A1 => gl_sig_green, A2 => gl_vgd_n_79, Z => G);
  gl_vgd_g1610 : AN2D4BWP7T port map(A1 => gl_sig_blue, A2 => gl_vgd_n_79, Z => B);
  gl_vgd_g1611 : INR4D0BWP7T port map(A1 => gl_vgd_n_71, B1 => gl_vgd_horizontal(1), B2 => gl_vgd_horizontal(0), B3 => gl_vgd_n_76, ZN => gl_sig_scale_h);
  gl_vgd_g1612 : AOI31D0BWP7T port map(A1 => gl_vgd_n_74, A2 => gl_vgd_horizontal(5), A3 => gl_vgd_horizontal(7), B => gl_vgd_n_78, ZN => gl_vgd_n_80);
  gl_vgd_g1613 : OR3D4BWP7T port map(A1 => gl_vgd_vertical(9), A2 => gl_vgd_n_69, A3 => gl_vgd_n_77, Z => V);
  gl_vgd_g1614 : IINR4D0BWP7T port map(A1 => gl_vgd_n_75, A2 => gl_vgd_n_69, B1 => gl_vgd_vertical(0), B2 => gl_vgd_vertical(9), ZN => gl_sig_scale_v);
  gl_vgd_g1615 : OAI31D0BWP7T port map(A1 => gl_vgd_horizontal(4), A2 => gl_vgd_horizontal(7), A3 => gl_vgd_n_72, B => gl_vgd_n_68, ZN => gl_vgd_n_78);
  gl_vgd_g1616 : INR3D0BWP7T port map(A1 => gl_vgd_n_69, B1 => gl_vgd_vertical(9), B2 => gl_vgd_n_76, ZN => gl_vgd_n_79);
  gl_vgd_g1617 : IND4D0BWP7T port map(A1 => gl_vgd_vertical(4), B1 => gl_vgd_vertical(3), B2 => gl_vgd_n_67, B3 => gl_vgd_n_70, ZN => gl_vgd_n_77);
  gl_vgd_g1618 : IND2D1BWP7T port map(A1 => gl_vgd_horizontal(9), B1 => gl_vgd_n_73, ZN => gl_vgd_n_76);
  gl_vgd_g1619 : NR3D0BWP7T port map(A1 => gl_vgd_n_67, A2 => gl_vgd_vertical(4), A3 => gl_vgd_vertical(3), ZN => gl_vgd_n_75);
  gl_vgd_g1620 : IOA21D1BWP7T port map(A1 => gl_vgd_horizontal(1), A2 => gl_vgd_horizontal(0), B => gl_vgd_n_71, ZN => gl_vgd_n_74);
  gl_vgd_g1621 : ND4D0BWP7T port map(A1 => gl_vgd_horizontal(5), A2 => gl_vgd_horizontal(7), A3 => gl_vgd_horizontal(8), A4 => gl_vgd_horizontal(6), ZN => gl_vgd_n_73);
  gl_vgd_g1622 : AO211D0BWP7T port map(A1 => gl_vgd_horizontal(2), A2 => gl_vgd_horizontal(1), B => gl_vgd_horizontal(5), C => gl_vgd_horizontal(3), Z => gl_vgd_n_72);
  gl_vgd_g1623 : MUX2ND0BWP7T port map(I0 => gl_vgd_vertical(1), I1 => gl_vgd_vertical(2), S => gl_vgd_vertical(0), ZN => gl_vgd_n_70);
  gl_vgd_g1624 : NR3D0BWP7T port map(A1 => gl_vgd_horizontal(4), A2 => gl_vgd_horizontal(2), A3 => gl_vgd_horizontal(3), ZN => gl_vgd_n_71);
  gl_vgd_g1625 : MAOI22D0BWP7T port map(A1 => gl_vgd_horizontal(7), A2 => gl_vgd_horizontal(6), B1 => gl_vgd_horizontal(7), B2 => gl_vgd_horizontal(6), ZN => gl_vgd_n_68);
  gl_vgd_g1626 : ND4D0BWP7T port map(A1 => gl_vgd_vertical(5), A2 => gl_vgd_vertical(7), A3 => gl_vgd_vertical(8), A4 => gl_vgd_vertical(6), ZN => gl_vgd_n_69);
  gl_vgd_g1627 : OR2D1BWP7T port map(A1 => gl_vgd_vertical(2), A2 => gl_vgd_vertical(1), Z => gl_vgd_n_67);
  gl_vgd_scale_horizontal_reg_8 : DFKCNQD1BWP7T port map(CP => clk, CN => gl_vgd_n_1, D => gl_vgd_horizontal_counter(8), Q => gl_vgd_horizontal(8));
  gl_vgd_vertical_reg_4 : DFKCNQD1BWP7T port map(CP => clk, CN => gl_vgd_n_1, D => gl_vgd_vertical_counter(4), Q => gl_vgd_vertical(4));
  gl_vgd_scale_horizontal_reg_3 : DFKCNQD1BWP7T port map(CP => clk, CN => gl_vgd_n_1, D => gl_vgd_horizontal_counter(3), Q => gl_vgd_horizontal(3));
  gl_vgd_vertical_reg_3 : DFKCNQD1BWP7T port map(CP => clk, CN => gl_vgd_n_1, D => gl_vgd_vertical_counter(3), Q => gl_vgd_vertical(3));
  gl_vgd_horizontal_reg_0 : DFKCNQD1BWP7T port map(CP => clk, CN => gl_vgd_n_1, D => gl_vgd_horizontal_counter(0), Q => gl_vgd_horizontal(0));
  gl_vgd_vertical_reg_2 : DFKCNQD1BWP7T port map(CP => clk, CN => gl_vgd_n_1, D => gl_vgd_vertical_counter(2), Q => gl_vgd_vertical(2));
  gl_vgd_vertical_reg_1 : DFKCNQD1BWP7T port map(CP => clk, CN => gl_vgd_n_1, D => gl_vgd_vertical_counter(1), Q => gl_vgd_vertical(1));
  gl_vgd_horizontal_reg_6 : DFKCNQD1BWP7T port map(CP => clk, CN => gl_vgd_n_1, D => gl_vgd_horizontal_counter(6), Q => gl_vgd_horizontal(6));
  gl_vgd_horizontal_reg_5 : DFKCNQD1BWP7T port map(CP => clk, CN => gl_vgd_n_1, D => gl_vgd_horizontal_counter(5), Q => gl_vgd_horizontal(5));
  gl_vgd_scale_horizontal_reg_1 : DFKCNQD1BWP7T port map(CP => clk, CN => gl_vgd_n_1, D => gl_vgd_horizontal_counter(1), Q => gl_vgd_horizontal(1));
  gl_vgd_scale_vertical_reg_7 : DFKCNQD1BWP7T port map(CP => clk, CN => gl_vgd_n_1, D => gl_vgd_vertical_counter(7), Q => gl_vgd_vertical(7));
  gl_vgd_scale_vertical_reg_8 : DFKCNQD1BWP7T port map(CP => clk, CN => gl_vgd_n_1, D => gl_vgd_vertical_counter(8), Q => gl_vgd_vertical(8));
  gl_vgd_scale_vertical_reg_6 : DFKCNQD1BWP7T port map(CP => clk, CN => gl_vgd_n_1, D => gl_vgd_vertical_counter(6), Q => gl_vgd_vertical(6));
  gl_vgd_vertical_reg_5 : DFKCNQD1BWP7T port map(CP => clk, CN => gl_vgd_n_1, D => gl_vgd_vertical_counter(5), Q => gl_vgd_vertical(5));
  gl_vgd_scale_horizontal_reg_4 : DFKCNQD1BWP7T port map(CP => clk, CN => gl_vgd_n_1, D => gl_vgd_horizontal_counter(4), Q => gl_vgd_horizontal(4));
  gl_vgd_horizontal_reg_9 : DFKCNQD1BWP7T port map(CP => clk, CN => gl_vgd_n_1, D => gl_vgd_horizontal_counter(9), Q => gl_vgd_horizontal(9));
  gl_vgd_scale_horizontal_reg_2 : DFKCNQD1BWP7T port map(CP => clk, CN => gl_vgd_n_1, D => gl_vgd_horizontal_counter(2), Q => gl_vgd_horizontal(2));
  gl_vgd_vertical_reg_0 : DFKCNQD1BWP7T port map(CP => clk, CN => gl_vgd_n_1, D => gl_vgd_vertical_counter(0), Q => gl_vgd_vertical(0));
  gl_vgd_scale_vertical_reg_9 : DFKCNQD1BWP7T port map(CP => clk, CN => gl_vgd_n_1, D => gl_vgd_vertical_counter(9), Q => gl_vgd_vertical(9));
  gl_vgd_horizontal_reg_7 : DFKCNQD1BWP7T port map(CP => clk, CN => gl_vgd_n_1, D => gl_vgd_horizontal_counter(7), Q => gl_vgd_horizontal(7));
  gl_vgd_g1648 : INVD1BWP7T port map(I => n_0, ZN => gl_vgd_n_1);
  gl_vgd_horizontal_counter_reg_0 : DFKCNQD1BWP7T port map(CP => clk, CN => gl_vgd_n_6, D => gl_vgd_n_41, Q => gl_vgd_horizontal_counter(0));
  gl_vgd_horizontal_counter_reg_1 : DFKCNQD1BWP7T port map(CP => clk, CN => gl_vgd_n_19, D => gl_vgd_n_41, Q => gl_vgd_horizontal_counter(1));
  gl_vgd_horizontal_counter_reg_2 : DFKCNQD1BWP7T port map(CP => clk, CN => gl_vgd_n_24, D => gl_vgd_n_41, Q => gl_vgd_horizontal_counter(2));
  gl_vgd_horizontal_counter_reg_3 : DFKCNQD1BWP7T port map(CP => clk, CN => gl_vgd_n_29, D => gl_vgd_n_41, Q => gl_vgd_horizontal_counter(3));
  gl_vgd_horizontal_counter_reg_4 : DFKCNQD1BWP7T port map(CP => clk, CN => gl_vgd_n_32, D => gl_vgd_n_41, Q => gl_vgd_horizontal_counter(4));
  gl_vgd_horizontal_counter_reg_5 : DFKCNQD1BWP7T port map(CP => clk, CN => gl_vgd_n_37, D => gl_vgd_n_41, Q => gl_vgd_horizontal_counter(5));
  gl_vgd_horizontal_counter_reg_6 : DFKCNQD1BWP7T port map(CP => clk, CN => gl_vgd_n_46, D => gl_vgd_n_41, Q => gl_vgd_horizontal_counter(6));
  gl_vgd_horizontal_counter_reg_7 : DFKCNQD1BWP7T port map(CP => clk, CN => gl_vgd_n_56, D => gl_vgd_n_41, Q => gl_vgd_horizontal_counter(7));
  gl_vgd_horizontal_counter_reg_8 : DFKCNQD1BWP7T port map(CP => clk, CN => gl_vgd_n_41, D => gl_vgd_n_62, Q => gl_vgd_horizontal_counter(8));
  gl_vgd_horizontal_counter_reg_9 : DFKCNQD1BWP7T port map(CP => clk, CN => gl_vgd_n_41, D => gl_vgd_n_65, Q => gl_vgd_horizontal_counter(9));
  gl_vgd_vertical_counter_reg_0 : DFXQD1BWP7T port map(CP => clk, DA => gl_vgd_n_44, DB => gl_vgd_n_43, SA => gl_vgd_vertical_counter(0), Q => gl_vgd_vertical_counter(0));
  gl_vgd_vertical_counter_reg_1 : DFQD1BWP7T port map(CP => clk, D => gl_vgd_n_51, Q => gl_vgd_vertical_counter(1));
  gl_vgd_vertical_counter_reg_2 : DFQD1BWP7T port map(CP => clk, D => gl_vgd_n_52, Q => gl_vgd_vertical_counter(2));
  gl_vgd_vertical_counter_reg_3 : DFQD1BWP7T port map(CP => clk, D => gl_vgd_n_49, Q => gl_vgd_vertical_counter(3));
  gl_vgd_vertical_counter_reg_4 : DFQD1BWP7T port map(CP => clk, D => gl_vgd_n_54, Q => gl_vgd_vertical_counter(4));
  gl_vgd_vertical_counter_reg_5 : DFQD1BWP7T port map(CP => clk, D => gl_vgd_n_53, Q => gl_vgd_vertical_counter(5));
  gl_vgd_vertical_counter_reg_6 : DFQD1BWP7T port map(CP => clk, D => gl_vgd_n_50, Q => gl_vgd_vertical_counter(6));
  gl_vgd_vertical_counter_reg_7 : DFQD1BWP7T port map(CP => clk, D => gl_vgd_n_57, Q => gl_vgd_vertical_counter(7));
  gl_vgd_vertical_counter_reg_9 : DFQD1BWP7T port map(CP => clk, D => gl_vgd_n_64, Q => gl_vgd_vertical_counter(9));
  gl_vgd_g1735 : MOAI22D0BWP7T port map(A1 => gl_vgd_n_63, A2 => gl_vgd_n_14, B1 => gl_vgd_n_63, B2 => gl_vgd_n_14, ZN => gl_vgd_n_65);
  gl_vgd_g1738 : AO22D0BWP7T port map(A1 => gl_vgd_n_58, A2 => gl_vgd_vertical_counter(9), B1 => gl_vgd_n_60, B2 => gl_vgd_n_43, Z => gl_vgd_n_64);
  gl_vgd_g1739 : HA1D0BWP7T port map(A => gl_vgd_n_11, B => gl_vgd_n_55, CO => gl_vgd_n_63, S => gl_vgd_n_62);
  gl_vgd_g1740 : AO21D0BWP7T port map(A1 => gl_vgd_n_58, A2 => gl_vgd_vertical_counter(8), B => gl_vgd_n_59, Z => gl_vgd_n_61);
  gl_vgd_g1742 : OAI31D0BWP7T port map(A1 => gl_vgd_vertical_counter(9), A2 => gl_vgd_n_2, A3 => gl_vgd_n_47, B => gl_vgd_n_15, ZN => gl_vgd_n_60);
  gl_vgd_g1744 : NR3D0BWP7T port map(A1 => gl_vgd_n_42, A2 => gl_vgd_n_47, A3 => gl_vgd_vertical_counter(8), ZN => gl_vgd_n_59);
  gl_vgd_g1745 : MOAI22D0BWP7T port map(A1 => gl_vgd_n_42, A2 => gl_vgd_n_48, B1 => gl_vgd_n_44, B2 => gl_vgd_vertical_counter(7), ZN => gl_vgd_n_57);
  gl_vgd_g1746 : AO21D0BWP7T port map(A1 => gl_vgd_n_43, A2 => gl_vgd_n_47, B => gl_vgd_n_44, Z => gl_vgd_n_58);
  gl_vgd_g1747 : HA1D0BWP7T port map(A => gl_vgd_n_13, B => gl_vgd_n_45, CO => gl_vgd_n_55, S => gl_vgd_n_56);
  gl_vgd_g1755 : MOAI22D0BWP7T port map(A1 => gl_vgd_n_42, A2 => gl_vgd_n_30, B1 => gl_vgd_n_44, B2 => gl_vgd_vertical_counter(4), ZN => gl_vgd_n_54);
  gl_vgd_g1756 : MOAI22D0BWP7T port map(A1 => gl_vgd_n_42, A2 => gl_vgd_n_34, B1 => gl_vgd_n_44, B2 => gl_vgd_vertical_counter(5), ZN => gl_vgd_n_53);
  gl_vgd_g1758 : MOAI22D0BWP7T port map(A1 => gl_vgd_n_42, A2 => gl_vgd_n_20, B1 => gl_vgd_n_44, B2 => gl_vgd_vertical_counter(2), ZN => gl_vgd_n_52);
  gl_vgd_g1759 : MOAI22D0BWP7T port map(A1 => gl_vgd_n_42, A2 => gl_vgd_n_0, B1 => gl_vgd_n_44, B2 => gl_vgd_vertical_counter(1), ZN => gl_vgd_n_51);
  gl_vgd_g1760 : MOAI22D0BWP7T port map(A1 => gl_vgd_n_42, A2 => gl_vgd_n_39, B1 => gl_vgd_n_44, B2 => gl_vgd_vertical_counter(6), ZN => gl_vgd_n_50);
  gl_vgd_g1761 : MOAI22D0BWP7T port map(A1 => gl_vgd_n_42, A2 => gl_vgd_n_25, B1 => gl_vgd_n_44, B2 => gl_vgd_vertical_counter(3), ZN => gl_vgd_n_49);
  gl_vgd_g1765 : MAOI22D0BWP7T port map(A1 => gl_vgd_n_38, A2 => gl_vgd_vertical_counter(7), B1 => gl_vgd_n_38, B2 => gl_vgd_vertical_counter(7), ZN => gl_vgd_n_48);
  gl_vgd_g1769 : HA1D0BWP7T port map(A => gl_vgd_n_12, B => gl_vgd_n_36, CO => gl_vgd_n_45, S => gl_vgd_n_46);
  gl_vgd_g1770 : IND2D1BWP7T port map(A1 => gl_vgd_n_38, B1 => gl_vgd_vertical_counter(7), ZN => gl_vgd_n_47);
  gl_vgd_g1771 : INVD1BWP7T port map(I => gl_vgd_n_43, ZN => gl_vgd_n_42);
  gl_vgd_g1772 : NR2D1BWP7T port map(A1 => gl_vgd_n_40, A2 => n_0, ZN => gl_vgd_n_44);
  gl_vgd_g1773 : NR2XD0BWP7T port map(A1 => gl_vgd_n_41, A2 => gl_vgd_n_26, ZN => gl_vgd_n_43);
  gl_vgd_g1774 : INVD1BWP7T port map(I => gl_vgd_n_41, ZN => gl_vgd_n_40);
  gl_vgd_g1775 : IND3D1BWP7T port map(A1 => gl_vgd_n_13, B1 => gl_vgd_n_11, B2 => gl_vgd_n_35, ZN => gl_vgd_n_41);
  gl_vgd_g1776 : MAOI22D0BWP7T port map(A1 => gl_vgd_n_31, A2 => gl_vgd_vertical_counter(6), B1 => gl_vgd_n_31, B2 => gl_vgd_vertical_counter(6), ZN => gl_vgd_n_39);
  gl_vgd_g1777 : HA1D0BWP7T port map(A => gl_vgd_n_8, B => gl_vgd_n_33, CO => gl_vgd_n_36, S => gl_vgd_n_37);
  gl_vgd_g1778 : IND2D1BWP7T port map(A1 => gl_vgd_n_31, B1 => gl_vgd_vertical_counter(6), ZN => gl_vgd_n_38);
  gl_vgd_g1779 : INR4D0BWP7T port map(A1 => gl_vgd_n_33, B1 => gl_vgd_n_14, B2 => gl_vgd_n_8, B3 => gl_vgd_n_12, ZN => gl_vgd_n_35);
  gl_vgd_g1780 : MAOI22D0BWP7T port map(A1 => gl_vgd_n_27, A2 => gl_vgd_vertical_counter(5), B1 => gl_vgd_n_27, B2 => gl_vgd_vertical_counter(5), ZN => gl_vgd_n_34);
  gl_vgd_g1781 : HA1D0BWP7T port map(A => gl_vgd_n_10, B => gl_vgd_n_28, CO => gl_vgd_n_33, S => gl_vgd_n_32);
  gl_vgd_g1782 : IND2D1BWP7T port map(A1 => gl_vgd_n_27, B1 => gl_vgd_vertical_counter(5), ZN => gl_vgd_n_31);
  gl_vgd_g1783 : MAOI22D0BWP7T port map(A1 => gl_vgd_n_22, A2 => gl_vgd_vertical_counter(4), B1 => gl_vgd_n_22, B2 => gl_vgd_vertical_counter(4), ZN => gl_vgd_n_30);
  gl_vgd_g1784 : HA1D0BWP7T port map(A => gl_vgd_n_4, B => gl_vgd_n_23, CO => gl_vgd_n_28, S => gl_vgd_n_29);
  gl_vgd_g1785 : IND2D1BWP7T port map(A1 => gl_vgd_n_22, B1 => gl_vgd_vertical_counter(4), ZN => gl_vgd_n_27);
  gl_vgd_g1786 : NR4D0BWP7T port map(A1 => gl_vgd_n_21, A2 => gl_vgd_vertical_counter(7), A3 => gl_vgd_vertical_counter(6), A4 => gl_vgd_vertical_counter(5), ZN => gl_vgd_n_26);
  gl_vgd_g1787 : MAOI22D0BWP7T port map(A1 => gl_vgd_n_17, A2 => gl_vgd_vertical_counter(3), B1 => gl_vgd_n_17, B2 => gl_vgd_vertical_counter(3), ZN => gl_vgd_n_25);
  gl_vgd_g1788 : HA1D0BWP7T port map(A => gl_vgd_n_3, B => gl_vgd_n_18, CO => gl_vgd_n_23, S => gl_vgd_n_24);
  gl_vgd_g1789 : IND2D1BWP7T port map(A1 => gl_vgd_n_17, B1 => gl_vgd_vertical_counter(3), ZN => gl_vgd_n_22);
  gl_vgd_g1790 : IND4D0BWP7T port map(A1 => gl_vgd_vertical_counter(4), B1 => gl_vgd_vertical_counter(2), B2 => gl_vgd_vertical_counter(3), B3 => gl_vgd_n_16, ZN => gl_vgd_n_21);
  gl_vgd_g1791 : MAOI22D0BWP7T port map(A1 => gl_vgd_n_9, A2 => gl_vgd_vertical_counter(2), B1 => gl_vgd_n_9, B2 => gl_vgd_vertical_counter(2), ZN => gl_vgd_n_20);
  gl_vgd_g1792 : HA1D0BWP7T port map(A => gl_vgd_n_7, B => gl_vgd_n_5, CO => gl_vgd_n_18, S => gl_vgd_n_19);
  gl_vgd_g1793 : IND2D1BWP7T port map(A1 => gl_vgd_n_9, B1 => gl_vgd_vertical_counter(2), ZN => gl_vgd_n_17);
  gl_vgd_g1794 : NR3D0BWP7T port map(A1 => gl_vgd_n_15, A2 => gl_vgd_vertical_counter(1), A3 => gl_vgd_vertical_counter(0), ZN => gl_vgd_n_16);
  gl_vgd_g1796 : ND2D1BWP7T port map(A1 => gl_vgd_n_2, A2 => gl_vgd_vertical_counter(9), ZN => gl_vgd_n_15);
  gl_vgd_g1797 : ND2D1BWP7T port map(A1 => gl_vgd_horizontal_counter(9), A2 => gl_vgd_n_1, ZN => gl_vgd_n_14);
  gl_vgd_g1798 : INR2XD0BWP7T port map(A1 => gl_vgd_horizontal_counter(4), B1 => n_0, ZN => gl_vgd_n_10);
  gl_vgd_g1799 : INR2D1BWP7T port map(A1 => gl_vgd_horizontal_counter(7), B1 => n_0, ZN => gl_vgd_n_13);
  gl_vgd_g1800 : INR2D1BWP7T port map(A1 => gl_vgd_horizontal_counter(6), B1 => n_0, ZN => gl_vgd_n_12);
  gl_vgd_g1801 : INR2D1BWP7T port map(A1 => gl_vgd_horizontal_counter(8), B1 => n_0, ZN => gl_vgd_n_11);
  gl_vgd_g1802 : INVD0BWP7T port map(I => gl_vgd_n_6, ZN => gl_vgd_n_7);
  gl_vgd_g1803 : CKAN2D1BWP7T port map(A1 => gl_vgd_horizontal_counter(1), A2 => gl_vgd_n_1, Z => gl_vgd_n_5);
  gl_vgd_g1804 : ND2D1BWP7T port map(A1 => gl_vgd_vertical_counter(1), A2 => gl_vgd_vertical_counter(0), ZN => gl_vgd_n_9);
  gl_vgd_g1805 : CKAN2D1BWP7T port map(A1 => gl_vgd_horizontal_counter(3), A2 => gl_vgd_n_1, Z => gl_vgd_n_4);
  gl_vgd_g1806 : CKAN2D1BWP7T port map(A1 => gl_vgd_horizontal_counter(2), A2 => gl_vgd_n_1, Z => gl_vgd_n_3);
  gl_vgd_g1807 : AN2D1BWP7T port map(A1 => gl_vgd_horizontal_counter(5), A2 => gl_vgd_n_1, Z => gl_vgd_n_8);
  gl_vgd_g1808 : ND2D1BWP7T port map(A1 => gl_vgd_horizontal_counter(0), A2 => gl_vgd_n_1, ZN => gl_vgd_n_6);
  gl_vgd_g2 : XNR2D1BWP7T port map(A1 => gl_vgd_vertical_counter(1), A2 => gl_vgd_vertical_counter(0), ZN => gl_vgd_n_0);
  gl_vgd_vertical_counter_reg_8 : DFD1BWP7T port map(CP => clk, D => gl_vgd_n_61, Q => gl_vgd_vertical_counter(8), QN => gl_vgd_n_2);
  ml_ms_mx2_g23 : MUX2D1BWP7T port map(I0 => ml_ms_cntReset25M_main, I1 => ml_ms_cntReset25M_send, S => ml_ms_mux_select_main, Z => ml_ms_cntReset25M);
  gl_gr_lg_y_grid_asked_reg_1 : LNQD1BWP7T port map(EN => gl_gr_lg_n_116, D => gl_gr_lg_n_115, Q => gl_sig_y(1));
  gl_gr_lg_y_grid_asked_reg_0 : LNQD1BWP7T port map(EN => gl_gr_lg_n_116, D => gl_gr_lg_n_114, Q => gl_sig_y(0));
  gl_gr_lg_x_grid_asked_reg_3 : LNQD1BWP7T port map(EN => gl_gr_lg_n_116, D => gl_gr_lg_n_110, Q => gl_sig_x(3));
  gl_gr_lg_x_grid_asked_reg_2 : LNQD1BWP7T port map(EN => gl_gr_lg_n_116, D => gl_gr_lg_n_111, Q => gl_sig_x(2));
  gl_gr_lg_x_grid_asked_reg_0 : LNQD1BWP7T port map(EN => gl_gr_lg_n_116, D => gl_gr_lg_n_113, Q => gl_sig_x(0));
  gl_gr_lg_x_grid_asked_reg_1 : LNQD1BWP7T port map(EN => gl_gr_lg_n_116, D => gl_gr_lg_n_107, Q => gl_sig_x(1));
  gl_gr_lg_y_grid_asked_reg_3 : LNQD1BWP7T port map(EN => gl_gr_lg_n_116, D => gl_gr_lg_n_108, Q => gl_sig_y(3));
  gl_gr_lg_y_grid_asked_reg_2 : LNQD1BWP7T port map(EN => gl_gr_lg_n_116, D => gl_gr_lg_n_112, Q => gl_sig_y(2));
  gl_gr_lg_g2072 : AO21D0BWP7T port map(A1 => gl_gr_lg_n_89, A2 => gl_gr_lg_n_155, B => gl_gr_lg_n_118, Z => gl_gr_lg_n_116);
  gl_gr_lg_g2073 : NR4D0BWP7T port map(A1 => gl_gr_lg_n_109, A2 => gl_gr_lg_n_85, A3 => gl_gr_lg_local_y(2), A4 => gl_gr_lg_local_y(3), ZN => gl_gr_lg_n_118);
  gl_gr_lg_g2074 : INR2D0BWP7T port map(A1 => gl_gr_lg_n_117, B1 => gl_gr_lg_n_85, ZN => gl_gr_lg_n_115);
  gl_gr_lg_g2075 : AN2D1BWP7T port map(A1 => gl_gr_lg_n_117, A2 => gl_gr_lg_local_y(0), Z => gl_gr_lg_n_114);
  gl_gr_lg_g2076 : INR2D0BWP7T port map(A1 => gl_gr_lg_n_117, B1 => gl_gr_lg_local_x(0), ZN => gl_gr_lg_n_113);
  gl_gr_lg_g2077 : INR2D0BWP7T port map(A1 => gl_gr_lg_n_117, B1 => gl_gr_lg_local_y(2), ZN => gl_gr_lg_n_112);
  gl_gr_lg_g2078 : OA21D0BWP7T port map(A1 => gl_gr_lg_n_99, A2 => gl_gr_lg_n_96, B => gl_gr_lg_n_117, Z => gl_gr_lg_n_111);
  gl_gr_lg_g2079 : NR3D0BWP7T port map(A1 => gl_gr_lg_n_106, A2 => gl_gr_lg_n_99, A3 => gl_gr_lg_n_1, ZN => gl_gr_lg_n_110);
  gl_gr_lg_g2080 : IND3D1BWP7T port map(A1 => gl_gr_lg_local_y(0), B1 => gl_gr_lg_n_102, B2 => gl_gr_lg_n_105, ZN => gl_gr_lg_n_109);
  gl_gr_lg_g2081 : INR2D0BWP7T port map(A1 => gl_gr_lg_n_117, B1 => gl_gr_lg_n_100, ZN => gl_gr_lg_n_108);
  gl_gr_lg_g2082 : OA21D0BWP7T port map(A1 => gl_gr_lg_n_90, A2 => gl_gr_lg_n_88, B => gl_gr_lg_n_117, Z => gl_gr_lg_n_107);
  gl_gr_lg_g2083 : NR4D0BWP7T port map(A1 => gl_gr_lg_n_104, A2 => gl_gr_lg_n_92, A3 => gl_gr_lg_n_95, A4 => gl_gr_lg_n_94, ZN => gl_gr_lg_n_155);
  gl_gr_lg_g2084 : INVD1BWP7T port map(I => gl_gr_lg_n_106, ZN => gl_gr_lg_n_117);
  gl_gr_lg_g2085 : OAI211D1BWP7T port map(A1 => gl_gr_lg_n_86, A2 => gl_gr_lg_n_100, B => gl_gr_lg_n_105, C => gl_gr_lg_n_101, ZN => gl_gr_lg_n_106);
  gl_gr_lg_g2086 : ND2D1BWP7T port map(A1 => gl_gr_lg_n_99, A2 => gl_gr_lg_n_1, ZN => gl_gr_lg_n_105);
  gl_gr_lg_g2087 : ND4D0BWP7T port map(A1 => gl_gr_lg_n_103, A2 => gl_gr_lg_n_98, A3 => gl_gr_lg_n_93, A4 => gl_gr_lg_n_97, ZN => gl_gr_lg_n_104);
  gl_gr_lg_g2088 : AOI211XD0BWP7T port map(A1 => gl_gr_lg_n_83, A2 => sig_logic_x(0), B => gl_gr_lg_n_91, C => gl_gr_lg_n_87, ZN => gl_gr_lg_n_103);
  gl_gr_lg_g2089 : ND4D0BWP7T port map(A1 => gl_gr_lg_n_83, A2 => gl_gr_lg_local_x(1), A3 => gl_gr_lg_local_x(2), A4 => gl_gr_lg_local_x(3), ZN => gl_gr_lg_n_102);
  gl_gr_lg_g2090 : OAI21D0BWP7T port map(A1 => gl_gr_lg_n_90, A2 => gl_gr_lg_local_x(2), B => gl_gr_lg_local_x(3), ZN => gl_gr_lg_n_101);
  gl_gr_lg_g2091 : XNR2D1BWP7T port map(A1 => gl_gr_lg_local_x(2), A2 => sig_logic_x(2), ZN => gl_gr_lg_n_98);
  gl_gr_lg_g2092 : MAOI22D0BWP7T port map(A1 => gl_gr_lg_n_1, A2 => sig_logic_x(3), B1 => gl_gr_lg_n_1, B2 => sig_logic_x(3), ZN => gl_gr_lg_n_97);
  gl_gr_lg_g2093 : INR2D0BWP7T port map(A1 => gl_gr_lg_local_x(2), B1 => gl_gr_lg_n_88, ZN => gl_gr_lg_n_96);
  gl_gr_lg_g2094 : CKXOR2D1BWP7T port map(A1 => gl_gr_lg_local_y(3), A2 => gl_gr_lg_local_y(2), Z => gl_gr_lg_n_100);
  gl_gr_lg_g2095 : INR2XD0BWP7T port map(A1 => gl_gr_lg_n_88, B1 => gl_gr_lg_local_x(2), ZN => gl_gr_lg_n_99);
  gl_gr_lg_g2096 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_n_85, A2 => sig_logic_y(1), B1 => gl_gr_lg_n_85, B2 => sig_logic_y(1), ZN => gl_gr_lg_n_95);
  gl_gr_lg_g2097 : CKXOR2D0BWP7T port map(A1 => gl_gr_lg_local_y(2), A2 => sig_logic_y(2), Z => gl_gr_lg_n_94);
  gl_gr_lg_g2098 : XNR2D1BWP7T port map(A1 => gl_gr_lg_local_x(1), A2 => sig_logic_x(1), ZN => gl_gr_lg_n_93);
  gl_gr_lg_g2099 : CKXOR2D0BWP7T port map(A1 => sig_logic_y(3), A2 => gl_gr_lg_local_y(3), Z => gl_gr_lg_n_92);
  gl_gr_lg_g2100 : CKXOR2D0BWP7T port map(A1 => gl_gr_lg_local_y(0), A2 => sig_logic_y(0), Z => gl_gr_lg_n_91);
  gl_gr_lg_g2101 : IND2D0BWP7T port map(A1 => gl_sig_rom(1), B1 => gl_sig_rom(0), ZN => gl_gr_lg_n_89);
  gl_gr_lg_g2102 : AN2D0BWP7T port map(A1 => gl_gr_lg_local_x(1), A2 => gl_gr_lg_local_x(0), Z => gl_gr_lg_n_90);
  gl_gr_lg_g2103 : NR2D0BWP7T port map(A1 => gl_gr_lg_n_83, A2 => sig_logic_x(0), ZN => gl_gr_lg_n_87);
  gl_gr_lg_g2104 : INR2D1BWP7T port map(A1 => gl_gr_lg_local_y(3), B1 => gl_gr_lg_local_y(1), ZN => gl_gr_lg_n_86);
  gl_gr_lg_g2105 : NR2XD0BWP7T port map(A1 => gl_gr_lg_local_x(1), A2 => gl_gr_lg_local_x(0), ZN => gl_gr_lg_n_88);
  gl_gr_lg_g2106 : INVD1BWP7T port map(I => gl_gr_lg_local_y(1), ZN => gl_gr_lg_n_85);
  gl_gr_lg_g2107 : INVD1BWP7T port map(I => gl_gr_lg_local_x(3), ZN => gl_gr_lg_n_1);
  gl_gr_lg_g2108 : INVD0BWP7T port map(I => gl_gr_lg_local_x(0), ZN => gl_gr_lg_n_83);
  gl_gr_lg_g2839 : IND4D0BWP7T port map(A1 => gl_gr_lg_n_81, B1 => gl_gr_lg_n_48, B2 => gl_gr_lg_n_26, B3 => gl_gr_lg_n_82, ZN => gl_sig_green);
  gl_gr_lg_g2840 : AOI211D1BWP7T port map(A1 => gl_gr_lg_n_56, A2 => gl_gr_lg_n_17, B => gl_gr_lg_n_80, C => gl_gr_lg_n_78, ZN => gl_gr_lg_n_82);
  gl_gr_lg_g2841 : OAI211D1BWP7T port map(A1 => gl_gr_lg_local_x(0), A2 => gl_gr_lg_n_65, B => gl_gr_lg_n_77, C => gl_gr_lg_n_74, ZN => gl_gr_lg_n_81);
  gl_gr_lg_g2842 : OAI31D0BWP7T port map(A1 => gl_gr_lg_countdown_case(6), A2 => gl_gr_lg_n_16, A3 => gl_gr_lg_n_51, B => gl_gr_lg_n_79, ZN => gl_gr_lg_n_80);
  gl_gr_lg_g2843 : AOI31D0BWP7T port map(A1 => gl_gr_lg_n_41, A2 => gl_gr_lg_n_54, A3 => gl_gr_lg_n_21, B => gl_gr_lg_n_76, ZN => gl_gr_lg_n_79);
  gl_gr_lg_g2844 : AO211D0BWP7T port map(A1 => gl_gr_lg_n_75, A2 => gl_gr_lg_n_0, B => gl_gr_lg_n_68, C => gl_gr_lg_n_73, Z => gl_gr_lg_n_78);
  gl_gr_lg_g2845 : AOI211D1BWP7T port map(A1 => gl_gr_lg_n_18, A2 => sig_output_color(1), B => gl_gr_lg_n_72, C => gl_gr_lg_n_58, ZN => gl_gr_lg_n_77);
  gl_gr_lg_g2846 : OAI222D0BWP7T port map(A1 => gl_gr_lg_n_71, A2 => gl_gr_lg_countdown_case(2), B1 => gl_gr_lg_local_x(0), B2 => gl_gr_lg_n_60, C1 => gl_gr_lg_n_44, C2 => gl_gr_lg_n_40, ZN => gl_gr_lg_n_76);
  gl_gr_lg_g2847 : OAI21D0BWP7T port map(A1 => gl_gr_lg_n_70, A2 => gl_gr_lg_countdown_case(8), B => gl_gr_lg_n_59, ZN => gl_gr_lg_n_75);
  gl_gr_lg_g2848 : AOI221D0BWP7T port map(A1 => gl_gr_lg_n_52, A2 => gl_gr_lg_n_36, B1 => gl_gr_lg_n_62, B2 => gl_gr_lg_n_7, C => gl_gr_lg_n_69, ZN => gl_gr_lg_n_74);
  gl_gr_lg_g2849 : OAI211D1BWP7T port map(A1 => gl_gr_lg_countdown_case(6), A2 => gl_gr_lg_n_55, B => gl_gr_lg_n_64, C => gl_gr_lg_n_67, ZN => gl_gr_lg_n_73);
  gl_gr_lg_g2850 : OAI33D1BWP7T port map(A1 => gl_gr_lg_local_x(0), A2 => gl_gr_lg_n_16, A3 => gl_gr_lg_n_63, B1 => gl_gr_lg_countdown_case(6), B2 => gl_gr_lg_n_31, B3 => gl_gr_lg_n_40, ZN => gl_gr_lg_n_72);
  gl_gr_lg_g2851 : IND3D1BWP7T port map(A1 => gl_gr_lg_countdown_case(1), B1 => gl_gr_lg_n_10, B2 => gl_gr_lg_n_66, ZN => gl_gr_lg_n_71);
  gl_gr_lg_g2852 : OAI21D0BWP7T port map(A1 => gl_gr_lg_n_21, A2 => gl_gr_lg_n_2, B => gl_gr_lg_n_66, ZN => gl_gr_lg_n_70);
  gl_gr_lg_g2853 : OAI33D1BWP7T port map(A1 => gl_gr_lg_countdown_case(5), A2 => gl_gr_lg_countdown_case(2), A3 => gl_gr_lg_n_53, B1 => gl_gr_lg_local_x(1), B2 => gl_gr_lg_n_20, B3 => gl_gr_lg_n_51, ZN => gl_gr_lg_n_69);
  gl_gr_lg_g2854 : OAI22D0BWP7T port map(A1 => gl_gr_lg_n_59, A2 => gl_gr_lg_local_x(0), B1 => gl_gr_lg_n_35, B2 => gl_gr_lg_n_45, ZN => gl_gr_lg_n_68);
  gl_gr_lg_g2855 : AOI22D0BWP7T port map(A1 => gl_gr_lg_n_43, A2 => gl_gr_lg_n_61, B1 => gl_gr_lg_n_41, B2 => gl_gr_lg_n_37, ZN => gl_gr_lg_n_67);
  gl_gr_lg_g2856 : OAI211D1BWP7T port map(A1 => gl_gr_lg_n_6, A2 => gl_gr_lg_n_3, B => gl_gr_lg_n_52, C => gl_gr_lg_n_1, ZN => gl_gr_lg_n_65);
  gl_gr_lg_g2857 : OAI31D0BWP7T port map(A1 => gl_gr_lg_local_x(0), A2 => gl_gr_lg_countdown_case(3), A3 => gl_gr_lg_n_47, B => gl_gr_lg_n_57, ZN => gl_gr_lg_n_66);
  gl_gr_lg_g2858 : OAI21D0BWP7T port map(A1 => gl_gr_lg_n_52, A2 => gl_gr_lg_n_156, B => gl_gr_lg_n_14, ZN => gl_gr_lg_n_64);
  gl_gr_lg_g2859 : OA21D0BWP7T port map(A1 => gl_gr_lg_n_49, A2 => gl_gr_lg_countdown_case(4), B => gl_gr_lg_n_51, Z => gl_gr_lg_n_63);
  gl_gr_lg_g2860 : OAI22D0BWP7T port map(A1 => gl_gr_lg_n_57, A2 => gl_gr_lg_n_9, B1 => gl_gr_lg_n_55, B2 => gl_gr_lg_countdown_case(5), ZN => gl_gr_lg_n_62);
  gl_gr_lg_g2861 : OAI31D0BWP7T port map(A1 => gl_gr_lg_countdown_case(3), A2 => gl_gr_lg_countdown_case(7), A3 => gl_gr_lg_n_25, B => gl_gr_lg_n_50, ZN => gl_gr_lg_n_61);
  gl_gr_lg_g2862 : IND3D1BWP7T port map(A1 => gl_gr_lg_n_51, B1 => gl_gr_lg_n_22, B2 => gl_gr_lg_n_28, ZN => gl_gr_lg_n_60);
  gl_gr_lg_g2863 : AOI21D0BWP7T port map(A1 => gl_gr_lg_countdown_case(8), A2 => gl_gr_lg_local_x(1), B => gl_gr_lg_n_55, ZN => gl_gr_lg_n_58);
  gl_gr_lg_g2864 : AOI21D0BWP7T port map(A1 => gl_gr_lg_n_43, A2 => gl_gr_lg_n_14, B => gl_gr_lg_n_56, ZN => gl_gr_lg_n_59);
  gl_gr_lg_g2865 : INVD0BWP7T port map(I => gl_gr_lg_n_56, ZN => gl_gr_lg_n_55);
  gl_gr_lg_g2866 : AO21D0BWP7T port map(A1 => gl_gr_lg_n_39, A2 => gl_gr_lg_n_7, B => gl_gr_lg_n_14, Z => gl_gr_lg_n_54);
  gl_gr_lg_g2867 : IND2D1BWP7T port map(A1 => gl_gr_lg_n_47, B1 => gl_gr_lg_n_38, ZN => gl_gr_lg_n_53);
  gl_gr_lg_g2868 : ND3D0BWP7T port map(A1 => gl_gr_lg_n_43, A2 => gl_gr_lg_n_17, A3 => gl_gr_lg_n_1, ZN => gl_gr_lg_n_57);
  gl_gr_lg_g2869 : NR2XD0BWP7T port map(A1 => gl_gr_lg_n_47, A2 => gl_gr_lg_countdown_case(9), ZN => gl_gr_lg_n_56);
  gl_gr_lg_g2870 : AOI33D1BWP7T port map(A1 => gl_gr_lg_n_29, A2 => gl_gr_lg_n_10, A3 => gl_gr_lg_n_6, B1 => gl_gr_lg_n_28, B2 => gl_gr_lg_n_13, B3 => gl_gr_lg_n_12, ZN => gl_gr_lg_n_50);
  gl_gr_lg_g2871 : AOI22D0BWP7T port map(A1 => gl_gr_lg_n_34, A2 => gl_gr_lg_n_38, B1 => gl_gr_lg_n_43, B2 => gl_gr_lg_n_12, ZN => gl_gr_lg_n_49);
  gl_gr_lg_g2872 : AOI22D0BWP7T port map(A1 => gl_gr_lg_n_41, A2 => gl_gr_lg_n_23, B1 => gl_gr_lg_n_24, B2 => gl_sig_ram(1), ZN => gl_gr_lg_n_48);
  gl_gr_lg_g2873 : OAI22D0BWP7T port map(A1 => gl_gr_lg_n_42, A2 => gl_gr_lg_countdown_case(8), B1 => gl_gr_lg_n_40, B2 => gl_gr_lg_countdown_case(7), ZN => gl_gr_lg_n_52);
  gl_gr_lg_g2874 : AOI21D0BWP7T port map(A1 => gl_gr_lg_n_43, A2 => gl_gr_lg_n_0, B => gl_gr_lg_n_41, ZN => gl_gr_lg_n_51);
  gl_gr_lg_g2875 : AO221D0BWP7T port map(A1 => gl_gr_lg_n_24, A2 => gl_sig_ram(0), B1 => gl_gr_lg_n_18, B2 => sig_output_color(0), C => gl_gr_lg_n_27, Z => gl_sig_red);
  gl_gr_lg_g2876 : AO221D0BWP7T port map(A1 => gl_gr_lg_n_24, A2 => gl_sig_ram(2), B1 => gl_gr_lg_n_18, B2 => sig_output_color(2), C => gl_gr_lg_n_27, Z => gl_sig_blue);
  gl_gr_lg_g2877 : IND2D1BWP7T port map(A1 => gl_gr_lg_countdown_case(10), B1 => gl_gr_lg_n_41, ZN => gl_gr_lg_n_47);
  gl_gr_lg_g2879 : OA22D0BWP7T port map(A1 => gl_gr_lg_n_30, A2 => gl_gr_lg_countdown_case(5), B1 => gl_gr_lg_local_x(3), B2 => gl_gr_lg_countdown_case(10), Z => gl_gr_lg_n_45);
  gl_gr_lg_g2880 : MAOI22D0BWP7T port map(A1 => gl_gr_lg_n_32, A2 => gl_gr_lg_n_22, B1 => gl_gr_lg_countdown_case(9), B2 => gl_gr_lg_local_x(3), ZN => gl_gr_lg_n_44);
  gl_gr_lg_g2881 : INVD0BWP7T port map(I => gl_gr_lg_n_43, ZN => gl_gr_lg_n_42);
  gl_gr_lg_g2882 : INVD1BWP7T port map(I => gl_gr_lg_n_41, ZN => gl_gr_lg_n_40);
  gl_gr_lg_g2883 : INR4D0BWP7T port map(A1 => gl_gr_lg_n_13, B1 => gl_gr_lg_local_x(3), B2 => gl_gr_lg_countdown_case(2), B3 => gl_gr_lg_countdown_case(4), ZN => gl_gr_lg_n_39);
  gl_gr_lg_g2884 : NR2XD0BWP7T port map(A1 => gl_gr_lg_n_35, A2 => gl_gr_lg_countdown_case(9), ZN => gl_gr_lg_n_43);
  gl_gr_lg_g2885 : NR2XD0BWP7T port map(A1 => gl_gr_lg_n_35, A2 => gl_gr_lg_local_x(2), ZN => gl_gr_lg_n_41);
  gl_gr_lg_g2886 : AOI211D1BWP7T port map(A1 => gl_gr_lg_n_15, A2 => gl_gr_lg_countdown_case(2), B => gl_gr_lg_n_25, C => gl_gr_lg_countdown_case(3), ZN => gl_gr_lg_n_37);
  gl_gr_lg_g2887 : OAI31D0BWP7T port map(A1 => gl_gr_lg_local_x(0), A2 => gl_gr_lg_local_x(1), A3 => gl_gr_lg_countdown_case(10), B => gl_gr_lg_n_33, ZN => gl_gr_lg_n_36);
  gl_gr_lg_g2888 : OAI32D1BWP7T port map(A1 => gl_gr_lg_countdown_case(3), A2 => gl_gr_lg_countdown_case(7), A3 => gl_gr_lg_n_9, B1 => gl_gr_lg_countdown_case(9), B2 => gl_gr_lg_n_15, ZN => gl_gr_lg_n_38);
  gl_gr_lg_g2889 : INVD0BWP7T port map(I => gl_gr_lg_n_35, ZN => gl_gr_lg_n_34);
  gl_gr_lg_g2890 : ND2D1BWP7T port map(A1 => gl_gr_lg_n_28, A2 => gl_gr_lg_n_17, ZN => gl_gr_lg_n_33);
  gl_gr_lg_g2891 : IOA21D1BWP7T port map(A1 => gl_gr_lg_n_8, A2 => gl_gr_lg_n_155, B => gl_gr_lg_n_118, ZN => gl_gr_lg_n_35);
  gl_gr_lg_g2892 : CKND1BWP7T port map(I => gl_gr_lg_n_31, ZN => gl_gr_lg_n_32);
  gl_gr_lg_g2893 : IND3D1BWP7T port map(A1 => gl_gr_lg_n_16, B1 => gl_gr_lg_n_10, B2 => gl_gr_lg_n_13, ZN => gl_gr_lg_n_30);
  gl_gr_lg_g2894 : AOI21D0BWP7T port map(A1 => gl_gr_lg_n_11, A2 => gl_gr_lg_countdown_case(1), B => gl_gr_lg_n_20, ZN => gl_gr_lg_n_29);
  gl_gr_lg_g2895 : AOI21D0BWP7T port map(A1 => gl_gr_lg_n_13, A2 => gl_gr_lg_n_19, B => gl_gr_lg_n_14, ZN => gl_gr_lg_n_31);
  gl_gr_lg_g2896 : CKND1BWP7T port map(I => gl_gr_lg_n_26, ZN => gl_gr_lg_n_27);
  gl_gr_lg_g2897 : NR2D1BWP7T port map(A1 => gl_gr_lg_n_9, A2 => gl_gr_lg_countdown_case(10), ZN => gl_gr_lg_n_28);
  gl_gr_lg_g2898 : ND2D1BWP7T port map(A1 => gl_gr_lg_n_18, A2 => gl_sig_rom(0), ZN => gl_gr_lg_n_26);
  gl_gr_lg_g2899 : AOI21D0BWP7T port map(A1 => gl_gr_lg_countdown_case(7), A2 => gl_gr_lg_local_x(1), B => gl_gr_lg_n_16, ZN => gl_gr_lg_n_23);
  gl_gr_lg_g2900 : IND2D1BWP7T port map(A1 => gl_gr_lg_n_16, B1 => gl_gr_lg_n_17, ZN => gl_gr_lg_n_25);
  gl_gr_lg_g2901 : OA21D0BWP7T port map(A1 => gl_sig_rom(0), A2 => gl_gr_lg_n_4, B => gl_gr_lg_n_117, Z => gl_gr_lg_n_24);
  gl_gr_lg_g2902 : CKND1BWP7T port map(I => gl_gr_lg_n_19, ZN => gl_gr_lg_n_20);
  gl_gr_lg_g2903 : CKND2D1BWP7T port map(A1 => gl_gr_lg_countdown_case(5), A2 => gl_gr_lg_countdown_case(4), ZN => gl_gr_lg_n_22);
  gl_gr_lg_g2904 : CKND2D1BWP7T port map(A1 => gl_gr_lg_countdown_case(1), A2 => gl_gr_lg_countdown_case(0), ZN => gl_gr_lg_n_21);
  gl_gr_lg_g2905 : NR2D1BWP7T port map(A1 => gl_gr_lg_countdown_case(8), A2 => gl_gr_lg_countdown_case(10), ZN => gl_gr_lg_n_19);
  gl_gr_lg_g2906 : CKAN2D1BWP7T port map(A1 => gl_sig_rom(1), A2 => gl_gr_lg_n_155, Z => gl_gr_lg_n_18);
  gl_gr_lg_g2907 : NR2XD0BWP7T port map(A1 => gl_gr_lg_countdown_case(4), A2 => gl_gr_lg_countdown_case(5), ZN => gl_gr_lg_n_17);
  gl_gr_lg_g2908 : OR2D1BWP7T port map(A1 => gl_gr_lg_countdown_case(8), A2 => gl_gr_lg_local_x(3), Z => gl_gr_lg_n_16);
  gl_gr_lg_g2909 : CKND1BWP7T port map(I => gl_gr_lg_n_12, ZN => gl_gr_lg_n_11);
  gl_gr_lg_g2910 : INVD1BWP7T port map(I => gl_gr_lg_n_10, ZN => gl_gr_lg_n_9);
  gl_gr_lg_g2912 : OR2D1BWP7T port map(A1 => gl_gr_lg_countdown_case(0), A2 => gl_gr_lg_countdown_case(1), Z => gl_gr_lg_n_15);
  gl_gr_lg_g2913 : NR2XD0BWP7T port map(A1 => gl_gr_lg_local_x(3), A2 => gl_gr_lg_local_x(1), ZN => gl_gr_lg_n_14);
  gl_gr_lg_g2914 : NR2D1BWP7T port map(A1 => gl_gr_lg_countdown_case(7), A2 => gl_gr_lg_local_x(0), ZN => gl_gr_lg_n_13);
  gl_gr_lg_g2915 : ND2D1BWP7T port map(A1 => gl_gr_lg_countdown_case(2), A2 => gl_gr_lg_countdown_case(3), ZN => gl_gr_lg_n_12);
  gl_gr_lg_g2916 : NR2D1BWP7T port map(A1 => gl_gr_lg_countdown_case(6), A2 => gl_gr_lg_local_x(1), ZN => gl_gr_lg_n_10);
  gl_gr_lg_g2917 : INVD0BWP7T port map(I => gl_gr_lg_countdown_case(3), ZN => gl_gr_lg_n_7);
  gl_gr_lg_g2918 : INVD0BWP7T port map(I => gl_gr_lg_countdown_case(5), ZN => gl_gr_lg_n_6);
  gl_gr_lg_g2920 : INVD0BWP7T port map(I => gl_gr_lg_n_155, ZN => gl_gr_lg_n_4);
  gl_gr_lg_g2921 : INVD0BWP7T port map(I => gl_gr_lg_countdown_case(6), ZN => gl_gr_lg_n_3);
  gl_gr_lg_g2922 : INVD0BWP7T port map(I => gl_gr_lg_countdown_case(2), ZN => gl_gr_lg_n_2);
  gl_gr_lg_g2924 : INVD0BWP7T port map(I => gl_gr_lg_countdown_case(7), ZN => gl_gr_lg_n_0);
  gl_gr_lg_g2925 : INVD0BWP7T port map(I => gl_sig_rom(0), ZN => gl_gr_lg_n_8);
  gl_gr_lg_g2 : INR2D1BWP7T port map(A1 => gl_gr_lg_n_12, B1 => gl_gr_lg_n_40, ZN => gl_gr_lg_n_156);
  gl_gr_lg_lcountdown_count_c_reg_7 : DFQD1BWP7T port map(CP => clk, D => gl_gr_lg_lcountdown_n_38, Q => gl_gr_lg_countdown_case(7));
  gl_gr_lg_lcountdown_g776 : OAI21D0BWP7T port map(A1 => gl_gr_lg_lcountdown_n_13, A2 => gl_gr_lg_lcountdown_n_36, B => gl_gr_lg_lcountdown_n_14, ZN => gl_gr_lg_lcountdown_n_38);
  gl_gr_lg_lcountdown_count_c_reg_6 : DFQD1BWP7T port map(CP => clk, D => gl_gr_lg_lcountdown_n_37, Q => gl_gr_lg_countdown_case(6));
  gl_gr_lg_lcountdown_count_c_reg_10 : DFQD1BWP7T port map(CP => clk, D => gl_gr_lg_lcountdown_n_35, Q => gl_gr_lg_countdown_case(10));
  gl_gr_lg_lcountdown_g779 : OAI21D0BWP7T port map(A1 => gl_gr_lg_lcountdown_n_13, A2 => gl_gr_lg_lcountdown_n_31, B => gl_gr_lg_lcountdown_n_14, ZN => gl_gr_lg_lcountdown_n_37);
  gl_gr_lg_lcountdown_g780 : MAOI22D0BWP7T port map(A1 => gl_gr_lg_lcountdown_n_30, A2 => gl_gr_lg_countdown_case(7), B1 => gl_gr_lg_lcountdown_n_30, B2 => gl_gr_lg_countdown_case(7), ZN => gl_gr_lg_lcountdown_n_36);
  gl_gr_lg_lcountdown_count_c_reg_9 : DFQD1BWP7T port map(CP => clk, D => gl_gr_lg_lcountdown_n_34, Q => gl_gr_lg_countdown_case(9));
  gl_gr_lg_lcountdown_g782 : OAI21D0BWP7T port map(A1 => gl_gr_lg_lcountdown_n_13, A2 => gl_gr_lg_lcountdown_n_33, B => gl_gr_lg_lcountdown_n_14, ZN => gl_gr_lg_lcountdown_n_35);
  gl_gr_lg_lcountdown_count_c_reg_5 : DFQD1BWP7T port map(CP => clk, D => gl_gr_lg_lcountdown_n_32, Q => gl_gr_lg_countdown_case(5));
  gl_gr_lg_lcountdown_g784 : OAI21D0BWP7T port map(A1 => gl_gr_lg_lcountdown_n_13, A2 => gl_gr_lg_lcountdown_n_28, B => gl_gr_lg_lcountdown_n_14, ZN => gl_gr_lg_lcountdown_n_34);
  gl_gr_lg_lcountdown_g785 : AOI21D0BWP7T port map(A1 => gl_gr_lg_lcountdown_n_23, A2 => gl_gr_lg_countdown_case(9), B => gl_gr_lg_countdown_case(10), ZN => gl_gr_lg_lcountdown_n_33);
  gl_gr_lg_lcountdown_g786 : OAI21D0BWP7T port map(A1 => gl_gr_lg_lcountdown_n_13, A2 => gl_gr_lg_lcountdown_n_26, B => gl_gr_lg_lcountdown_n_14, ZN => gl_gr_lg_lcountdown_n_32);
  gl_gr_lg_lcountdown_g787 : MAOI22D0BWP7T port map(A1 => gl_gr_lg_lcountdown_n_25, A2 => gl_gr_lg_countdown_case(6), B1 => gl_gr_lg_lcountdown_n_25, B2 => gl_gr_lg_countdown_case(6), ZN => gl_gr_lg_lcountdown_n_31);
  gl_gr_lg_lcountdown_count_c_reg_8 : DFQD1BWP7T port map(CP => clk, D => gl_gr_lg_lcountdown_n_29, Q => gl_gr_lg_countdown_case(8));
  gl_gr_lg_lcountdown_g789 : IND2D1BWP7T port map(A1 => gl_gr_lg_lcountdown_n_25, B1 => gl_gr_lg_countdown_case(6), ZN => gl_gr_lg_lcountdown_n_30);
  gl_gr_lg_lcountdown_count_c_reg_4 : DFQD1BWP7T port map(CP => clk, D => gl_gr_lg_lcountdown_n_27, Q => gl_gr_lg_countdown_case(4));
  gl_gr_lg_lcountdown_g791 : OAI21D0BWP7T port map(A1 => gl_gr_lg_lcountdown_n_13, A2 => gl_gr_lg_lcountdown_n_24, B => gl_gr_lg_lcountdown_n_14, ZN => gl_gr_lg_lcountdown_n_29);
  gl_gr_lg_lcountdown_g792 : XNR2D1BWP7T port map(A1 => gl_gr_lg_lcountdown_n_23, A2 => gl_gr_lg_countdown_case(9), ZN => gl_gr_lg_lcountdown_n_28);
  gl_gr_lg_lcountdown_g793 : OAI21D0BWP7T port map(A1 => gl_gr_lg_lcountdown_n_13, A2 => gl_gr_lg_lcountdown_n_21, B => gl_gr_lg_lcountdown_n_14, ZN => gl_gr_lg_lcountdown_n_27);
  gl_gr_lg_lcountdown_g794 : MAOI22D0BWP7T port map(A1 => gl_gr_lg_lcountdown_n_19, A2 => gl_gr_lg_countdown_case(5), B1 => gl_gr_lg_lcountdown_n_19, B2 => gl_gr_lg_countdown_case(5), ZN => gl_gr_lg_lcountdown_n_26);
  gl_gr_lg_lcountdown_g795 : IND2D1BWP7T port map(A1 => gl_gr_lg_lcountdown_n_19, B1 => gl_gr_lg_countdown_case(5), ZN => gl_gr_lg_lcountdown_n_25);
  gl_gr_lg_lcountdown_count_c_reg_3 : DFQD1BWP7T port map(CP => clk, D => gl_gr_lg_lcountdown_n_22, Q => gl_gr_lg_countdown_case(3));
  gl_gr_lg_lcountdown_g797 : MAOI22D0BWP7T port map(A1 => gl_gr_lg_lcountdown_n_20, A2 => gl_gr_lg_countdown_case(8), B1 => gl_gr_lg_lcountdown_n_20, B2 => gl_gr_lg_countdown_case(8), ZN => gl_gr_lg_lcountdown_n_24);
  gl_gr_lg_lcountdown_count_c_reg_1 : DFQD1BWP7T port map(CP => clk, D => gl_gr_lg_lcountdown_n_18, Q => gl_gr_lg_countdown_case(1));
  gl_gr_lg_lcountdown_count_c_reg_2 : DFQD1BWP7T port map(CP => clk, D => gl_gr_lg_lcountdown_n_16, Q => gl_gr_lg_countdown_case(2));
  gl_gr_lg_lcountdown_count_c_reg_0 : DFQD1BWP7T port map(CP => clk, D => gl_gr_lg_lcountdown_n_17, Q => gl_gr_lg_countdown_case(0));
  gl_gr_lg_lcountdown_g801 : OAI21D0BWP7T port map(A1 => gl_gr_lg_lcountdown_n_13, A2 => gl_gr_lg_lcountdown_n_12, B => gl_gr_lg_lcountdown_n_14, ZN => gl_gr_lg_lcountdown_n_22);
  gl_gr_lg_lcountdown_g802 : MAOI22D0BWP7T port map(A1 => gl_gr_lg_lcountdown_n_11, A2 => gl_gr_lg_countdown_case(4), B1 => gl_gr_lg_lcountdown_n_11, B2 => gl_gr_lg_countdown_case(4), ZN => gl_gr_lg_lcountdown_n_21);
  gl_gr_lg_lcountdown_g803 : INR2XD0BWP7T port map(A1 => gl_gr_lg_countdown_case(8), B1 => gl_gr_lg_lcountdown_n_20, ZN => gl_gr_lg_lcountdown_n_23);
  gl_gr_lg_lcountdown_countdown_aan_reg : DFQD1BWP7T port map(CP => clk, D => gl_gr_lg_lcountdown_n_15, Q => gl_sig_countdown_aan);
  gl_gr_lg_lcountdown_g805 : OR2D1BWP7T port map(A1 => gl_gr_lg_lcountdown_n_11, A2 => gl_gr_lg_lcountdown_n_3, Z => gl_gr_lg_lcountdown_n_20);
  gl_gr_lg_lcountdown_g806 : IND2D1BWP7T port map(A1 => gl_gr_lg_lcountdown_n_11, B1 => gl_gr_lg_countdown_case(4), ZN => gl_gr_lg_lcountdown_n_19);
  gl_gr_lg_lcountdown_g807 : OAI21D0BWP7T port map(A1 => gl_gr_lg_lcountdown_n_13, A2 => gl_gr_lg_lcountdown_n_6, B => gl_gr_lg_lcountdown_n_14, ZN => gl_gr_lg_lcountdown_n_18);
  gl_gr_lg_lcountdown_g808 : OAI21D0BWP7T port map(A1 => gl_gr_lg_lcountdown_n_13, A2 => gl_gr_lg_lcountdown_n_2, B => gl_gr_lg_lcountdown_n_14, ZN => gl_gr_lg_lcountdown_n_17);
  gl_gr_lg_lcountdown_g809 : OAI21D0BWP7T port map(A1 => gl_gr_lg_lcountdown_n_13, A2 => gl_gr_lg_lcountdown_n_9, B => gl_gr_lg_lcountdown_n_14, ZN => gl_gr_lg_lcountdown_n_16);
  gl_gr_lg_lcountdown_g810 : IOA21D1BWP7T port map(A1 => gl_gr_lg_lcountdown_n_1, A2 => gl_sig_countdown_aan, B => gl_gr_lg_lcountdown_n_13, ZN => gl_gr_lg_lcountdown_n_15);
  gl_gr_lg_lcountdown_g811 : IND3D1BWP7T port map(A1 => gl_gr_lg_lcountdown_n_1, B1 => gl_gr_lg_countdown_case(9), B2 => gl_gr_lg_lcountdown_n_10, ZN => gl_gr_lg_lcountdown_n_14);
  gl_gr_lg_lcountdown_g812 : MAOI22D0BWP7T port map(A1 => gl_gr_lg_lcountdown_n_8, A2 => gl_gr_lg_countdown_case(3), B1 => gl_gr_lg_lcountdown_n_8, B2 => gl_gr_lg_countdown_case(3), ZN => gl_gr_lg_lcountdown_n_12);
  gl_gr_lg_lcountdown_g813 : AO21D0BWP7T port map(A1 => gl_gr_lg_lcountdown_n_10, A2 => gl_gr_lg_countdown_case(9), B => gl_gr_lg_lcountdown_n_1, Z => gl_gr_lg_lcountdown_n_13);
  gl_gr_lg_lcountdown_g814 : IND2D1BWP7T port map(A1 => gl_gr_lg_lcountdown_n_8, B1 => gl_gr_lg_countdown_case(3), ZN => gl_gr_lg_lcountdown_n_11);
  gl_gr_lg_lcountdown_g815 : AN4D1BWP7T port map(A1 => gl_gr_lg_lcountdown_n_7, A2 => gl_gr_lg_countdown_case(2), A3 => gl_gr_lg_countdown_case(3), A4 => gl_gr_lg_countdown_case(8), Z => gl_gr_lg_lcountdown_n_10);
  gl_gr_lg_lcountdown_g816 : MAOI22D0BWP7T port map(A1 => gl_gr_lg_lcountdown_n_5, A2 => gl_gr_lg_countdown_case(2), B1 => gl_gr_lg_lcountdown_n_5, B2 => gl_gr_lg_countdown_case(2), ZN => gl_gr_lg_lcountdown_n_9);
  gl_gr_lg_lcountdown_g817 : IND2D1BWP7T port map(A1 => gl_gr_lg_lcountdown_n_5, B1 => gl_gr_lg_countdown_case(2), ZN => gl_gr_lg_lcountdown_n_8);
  gl_gr_lg_lcountdown_g818 : AN4D0BWP7T port map(A1 => gl_gr_lg_lcountdown_n_4, A2 => gl_gr_lg_countdown_case(10), A3 => gl_gr_lg_countdown_case(0), A4 => gl_gr_lg_countdown_case(1), Z => gl_gr_lg_lcountdown_n_7);
  gl_gr_lg_lcountdown_g819 : MAOI22D0BWP7T port map(A1 => gl_gr_lg_lcountdown_n_0, A2 => gl_gr_lg_countdown_case(1), B1 => gl_gr_lg_lcountdown_n_0, B2 => gl_gr_lg_countdown_case(1), ZN => gl_gr_lg_lcountdown_n_6);
  gl_gr_lg_lcountdown_g820 : IND2D1BWP7T port map(A1 => gl_gr_lg_lcountdown_n_0, B1 => gl_gr_lg_countdown_case(1), ZN => gl_gr_lg_lcountdown_n_5);
  gl_gr_lg_lcountdown_g821 : CKND1BWP7T port map(I => gl_gr_lg_lcountdown_n_3, ZN => gl_gr_lg_lcountdown_n_4);
  gl_gr_lg_lcountdown_g822 : ND4D0BWP7T port map(A1 => gl_gr_lg_countdown_case(6), A2 => gl_gr_lg_countdown_case(5), A3 => gl_gr_lg_countdown_case(7), A4 => gl_gr_lg_countdown_case(4), ZN => gl_gr_lg_lcountdown_n_3);
  gl_gr_lg_lcountdown_g823 : XNR2D1BWP7T port map(A1 => gl_gr_lg_countdown_case(0), A2 => gl_gr_lg_lcountdown_sig_edge_fall, ZN => gl_gr_lg_lcountdown_n_2);
  gl_gr_lg_lcountdown_g824 : OR2D1BWP7T port map(A1 => sig_middelsteknop, A2 => n_0, Z => gl_gr_lg_lcountdown_n_1);
  gl_gr_lg_lcountdown_g825 : ND2D1BWP7T port map(A1 => gl_gr_lg_countdown_case(0), A2 => gl_gr_lg_lcountdown_sig_edge_fall, ZN => gl_gr_lg_lcountdown_n_0);
  gl_gr_lg_lcountdown_l_edge_g12 : NR2XD0BWP7T port map(A1 => gl_gr_lg_lcountdown_l_edge_reg2, A2 => gl_gr_lg_lcountdown_l_edge_reg1, ZN => gl_gr_lg_lcountdown_sig_edge_fall);
  gl_gr_lg_lcountdown_l_edge_reg2_reg : DFD0BWP7T port map(CP => clk, D => gl_gr_lg_lcountdown_l_edge_reg1, Q => UNCONNECTED1, QN => gl_gr_lg_lcountdown_l_edge_reg2);
  gl_gr_lg_lcountdown_l_edge_reg1_reg : DFQD1BWP7T port map(CP => clk, D => V, Q => gl_gr_lg_lcountdown_l_edge_reg1);
  gl_gr_lg_le_g165 : INVD0BWP7T port map(I => gl_gr_lg_le_n_42, ZN => gl_gr_lg_le_n_41);
  gl_gr_lg_le_g366 : AN4D1BWP7T port map(A1 => gl_gr_lg_le_n_40, A2 => gl_gr_lg_le_n_39, A3 => gl_gr_lg_le_n_37, A4 => gl_gr_lg_le_n_32, Z => gl_gr_lg_le_n_42);
  gl_gr_lg_le_g367 : NR4D0BWP7T port map(A1 => gl_gr_lg_le_n_31, A2 => gl_gr_lg_le_n_33, A3 => gl_gr_lg_le_n_38, A4 => gl_gr_lg_le_n_36, ZN => gl_gr_lg_le_n_40);
  gl_gr_lg_le_g368 : NR2XD0BWP7T port map(A1 => gl_gr_lg_le_n_34, A2 => gl_gr_lg_le_n_35, ZN => gl_gr_lg_le_n_39);
  gl_gr_lg_le_g369 : CKXOR2D0BWP7T port map(A1 => sig_logic_y(1), A2 => gl_gr_lg_local_y(1), Z => gl_gr_lg_le_n_38);
  gl_gr_lg_le_g370 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_local_x(3), A2 => sig_logic_x(3), B1 => gl_gr_lg_local_x(3), B2 => sig_logic_x(3), ZN => gl_gr_lg_le_n_37);
  gl_gr_lg_le_g371 : CKXOR2D0BWP7T port map(A1 => sig_logic_y(2), A2 => gl_gr_lg_local_y(2), Z => gl_gr_lg_le_n_36);
  gl_gr_lg_le_g372 : MAOI22D0BWP7T port map(A1 => sig_logic_x(2), A2 => gl_gr_lg_local_x(2), B1 => sig_logic_x(2), B2 => gl_gr_lg_local_x(2), ZN => gl_gr_lg_le_n_35);
  gl_gr_lg_le_g373 : MAOI22D0BWP7T port map(A1 => gl_gr_lg_local_x(1), A2 => sig_logic_x(1), B1 => gl_gr_lg_local_x(1), B2 => sig_logic_x(1), ZN => gl_gr_lg_le_n_34);
  gl_gr_lg_le_g374 : CKXOR2D0BWP7T port map(A1 => sig_logic_y(0), A2 => gl_gr_lg_local_y(0), Z => gl_gr_lg_le_n_33);
  gl_gr_lg_le_g375 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_local_x(0), A2 => sig_logic_x(0), B1 => gl_gr_lg_local_x(0), B2 => sig_logic_x(0), ZN => gl_gr_lg_le_n_32);
  gl_gr_lg_le_g376 : CKXOR2D0BWP7T port map(A1 => sig_logic_y(3), A2 => gl_gr_lg_local_y(3), Z => gl_gr_lg_le_n_31);
  gl_gr_lg_le_new_count_e_reg_9 : LNQD1BWP7T port map(EN => gl_gr_lg_le_n_29, D => gl_gr_lg_le_n_30, Q => gl_gr_lg_le_new_count_e(9));
  gl_gr_lg_le_g464 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_le_n_27, A2 => gl_sig_e(9), B1 => gl_gr_lg_le_n_27, B2 => gl_sig_e(9), ZN => gl_gr_lg_le_n_30);
  gl_gr_lg_le_new_count_e_reg_8 : LNQD1BWP7T port map(EN => gl_gr_lg_le_n_29, D => gl_gr_lg_le_n_28, Q => gl_gr_lg_le_new_count_e(8));
  gl_gr_lg_le_g466 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_le_n_25, A2 => gl_sig_e(8), B1 => gl_gr_lg_le_n_25, B2 => gl_sig_e(8), ZN => gl_gr_lg_le_n_28);
  gl_gr_lg_le_new_count_e_reg_7 : LNQD1BWP7T port map(EN => gl_gr_lg_le_n_29, D => gl_gr_lg_le_n_26, Q => gl_gr_lg_le_new_count_e(7));
  gl_gr_lg_le_g468 : IND2D1BWP7T port map(A1 => gl_gr_lg_le_n_25, B1 => gl_sig_e(8), ZN => gl_gr_lg_le_n_27);
  gl_gr_lg_le_g469 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_le_n_23, A2 => gl_sig_e(7), B1 => gl_gr_lg_le_n_23, B2 => gl_sig_e(7), ZN => gl_gr_lg_le_n_26);
  gl_gr_lg_le_new_count_e_reg_6 : LNQD1BWP7T port map(EN => gl_gr_lg_le_n_29, D => gl_gr_lg_le_n_24, Q => gl_gr_lg_le_new_count_e(6));
  gl_gr_lg_le_g471 : IND2D1BWP7T port map(A1 => gl_gr_lg_le_n_23, B1 => gl_sig_e(7), ZN => gl_gr_lg_le_n_25);
  gl_gr_lg_le_g472 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_le_n_21, A2 => gl_sig_e(6), B1 => gl_gr_lg_le_n_21, B2 => gl_sig_e(6), ZN => gl_gr_lg_le_n_24);
  gl_gr_lg_le_new_count_e_reg_5 : LNQD1BWP7T port map(EN => gl_gr_lg_le_n_29, D => gl_gr_lg_le_n_22, Q => gl_gr_lg_le_new_count_e(5));
  gl_gr_lg_le_g474 : IND2D1BWP7T port map(A1 => gl_gr_lg_le_n_21, B1 => gl_sig_e(6), ZN => gl_gr_lg_le_n_23);
  gl_gr_lg_le_g475 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_le_n_19, A2 => gl_sig_e(5), B1 => gl_gr_lg_le_n_19, B2 => gl_sig_e(5), ZN => gl_gr_lg_le_n_22);
  gl_gr_lg_le_new_count_e_reg_4 : LNQD1BWP7T port map(EN => gl_gr_lg_le_n_29, D => gl_gr_lg_le_n_20, Q => gl_gr_lg_le_new_count_e(4));
  gl_gr_lg_le_g477 : IND2D1BWP7T port map(A1 => gl_gr_lg_le_n_19, B1 => gl_sig_e(5), ZN => gl_gr_lg_le_n_21);
  gl_gr_lg_le_g478 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_le_n_17, A2 => gl_sig_e(4), B1 => gl_gr_lg_le_n_17, B2 => gl_sig_e(4), ZN => gl_gr_lg_le_n_20);
  gl_gr_lg_le_new_count_e_reg_3 : LNQD1BWP7T port map(EN => gl_gr_lg_le_n_29, D => gl_gr_lg_le_n_18, Q => gl_gr_lg_le_new_count_e(3));
  gl_gr_lg_le_g480 : IND2D1BWP7T port map(A1 => gl_gr_lg_le_n_17, B1 => gl_sig_e(4), ZN => gl_gr_lg_le_n_19);
  gl_gr_lg_le_g481 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_le_n_15, A2 => gl_sig_e(3), B1 => gl_gr_lg_le_n_15, B2 => gl_sig_e(3), ZN => gl_gr_lg_le_n_18);
  gl_gr_lg_le_new_count_e_reg_2 : LNQD1BWP7T port map(EN => gl_gr_lg_le_n_29, D => gl_gr_lg_le_n_16, Q => gl_gr_lg_le_new_count_e(2));
  gl_gr_lg_le_g483 : IND2D1BWP7T port map(A1 => gl_gr_lg_le_n_15, B1 => gl_sig_e(3), ZN => gl_gr_lg_le_n_17);
  gl_gr_lg_le_g484 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_le_n_13, A2 => gl_sig_e(2), B1 => gl_gr_lg_le_n_13, B2 => gl_sig_e(2), ZN => gl_gr_lg_le_n_16);
  gl_gr_lg_le_new_count_e_reg_1 : LNQD1BWP7T port map(EN => gl_gr_lg_le_n_29, D => gl_gr_lg_le_n_14, Q => gl_gr_lg_le_new_count_e(1));
  gl_gr_lg_le_g486 : IND2D1BWP7T port map(A1 => gl_gr_lg_le_n_13, B1 => gl_sig_e(2), ZN => gl_gr_lg_le_n_15);
  gl_gr_lg_le_g487 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_le_n_11, A2 => gl_sig_e(1), B1 => gl_gr_lg_le_n_11, B2 => gl_sig_e(1), ZN => gl_gr_lg_le_n_14);
  gl_gr_lg_le_new_count_e_reg_0 : LNQD1BWP7T port map(EN => gl_gr_lg_le_n_29, D => gl_gr_lg_le_n_12, Q => gl_gr_lg_le_new_count_e(0));
  gl_gr_lg_le_g489 : IND2D1BWP7T port map(A1 => gl_gr_lg_le_n_11, B1 => gl_sig_e(1), ZN => gl_gr_lg_le_n_13);
  gl_gr_lg_le_g490 : AOI21D0BWP7T port map(A1 => clk, A2 => gl_gr_lg_le_n_42, B => gl_gr_lg_le_n_41, ZN => gl_gr_lg_le_n_29);
  gl_gr_lg_le_g491 : CKXOR2D1BWP7T port map(A1 => gl_gr_lg_le_n_42, A2 => gl_sig_e(0), Z => gl_gr_lg_le_n_12);
  gl_gr_lg_le_g492 : ND2D1BWP7T port map(A1 => gl_gr_lg_le_n_42, A2 => gl_sig_e(0), ZN => gl_gr_lg_le_n_11);
  gl_gr_lg_le_count_e_reg_2 : DFKCNQD2BWP7T port map(CP => clk, CN => gl_gr_lg_le_new_count_e(2), D => gl_gr_lg_le_n_10, Q => gl_sig_e(2));
  gl_gr_lg_le_count_e_reg_1 : DFKCNQD2BWP7T port map(CP => clk, CN => gl_gr_lg_le_new_count_e(1), D => gl_gr_lg_le_n_10, Q => gl_sig_e(1));
  gl_gr_lg_le_count_e_reg_0 : DFKCNQD2BWP7T port map(CP => clk, CN => gl_gr_lg_le_new_count_e(0), D => gl_gr_lg_le_n_10, Q => gl_sig_e(0));
  gl_gr_lg_le_count_e_reg_3 : DFKCNQD1BWP7T port map(CP => clk, CN => gl_gr_lg_le_new_count_e(3), D => gl_gr_lg_le_n_10, Q => gl_sig_e(3));
  gl_gr_lg_le_count_e_reg_4 : DFKCNQD1BWP7T port map(CP => clk, CN => gl_gr_lg_le_n_10, D => gl_gr_lg_le_new_count_e(4), Q => gl_sig_e(4));
  gl_gr_lg_le_count_e_reg_7 : DFKCNQD1BWP7T port map(CP => clk, CN => gl_gr_lg_le_n_10, D => gl_gr_lg_le_new_count_e(7), Q => gl_sig_e(7));
  gl_gr_lg_le_count_e_reg_6 : DFKCNQD1BWP7T port map(CP => clk, CN => gl_gr_lg_le_n_10, D => gl_gr_lg_le_new_count_e(6), Q => gl_sig_e(6));
  gl_gr_lg_le_count_e_reg_5 : DFKCNQD1BWP7T port map(CP => clk, CN => gl_gr_lg_le_n_10, D => gl_gr_lg_le_new_count_e(5), Q => gl_sig_e(5));
  gl_gr_lg_le_count_e_reg_8 : DFKCNQD1BWP7T port map(CP => clk, CN => gl_gr_lg_le_n_10, D => gl_gr_lg_le_new_count_e(8), Q => gl_sig_e(8));
  gl_gr_lg_le_count_e_reg_9 : DFKCNQD1BWP7T port map(CP => clk, CN => gl_gr_lg_le_n_10, D => gl_gr_lg_le_new_count_e(9), Q => gl_sig_e(9));
  gl_gr_lg_le_g432 : NR4D0BWP7T port map(A1 => gl_gr_lg_le_n_9, A2 => gl_gr_lg_le_n_6, A3 => gl_gr_lg_le_n_4, A4 => n_0, ZN => gl_gr_lg_le_n_10);
  gl_gr_lg_le_g433 : ND4D0BWP7T port map(A1 => gl_gr_lg_le_n_8, A2 => gl_gr_lg_le_n_3, A3 => gl_gr_lg_le_n_2, A4 => gl_gr_lg_le_n_1, ZN => gl_gr_lg_le_n_9);
  gl_gr_lg_le_g434 : NR3D0BWP7T port map(A1 => gl_gr_lg_le_n_0, A2 => gl_gr_lg_le_n_5, A3 => gl_gr_lg_le_n_7, ZN => gl_gr_lg_le_n_8);
  gl_gr_lg_le_x_old_reg_2 : DFXQD1BWP7T port map(CP => clk, DA => gl_gr_lg_le_x_old(2), DB => sig_logic_x(2), SA => n_0, Q => gl_gr_lg_le_x_old(2));
  gl_gr_lg_le_x_old_reg_1 : DFXQD1BWP7T port map(CP => clk, DA => gl_gr_lg_le_x_old(1), DB => sig_logic_x(1), SA => n_0, Q => gl_gr_lg_le_x_old(1));
  gl_gr_lg_le_x_old_reg_0 : DFXQD1BWP7T port map(CP => clk, DA => gl_gr_lg_le_x_old(0), DB => sig_logic_x(0), SA => n_0, Q => gl_gr_lg_le_x_old(0));
  gl_gr_lg_le_x_old_reg_3 : DFXQD1BWP7T port map(CP => clk, DA => gl_gr_lg_le_x_old(3), DB => sig_logic_x(3), SA => n_0, Q => gl_gr_lg_le_x_old(3));
  gl_gr_lg_le_y_old_reg_2 : DFXQD1BWP7T port map(CP => clk, DA => gl_gr_lg_le_y_old(2), DB => sig_logic_y(2), SA => n_0, Q => gl_gr_lg_le_y_old(2));
  gl_gr_lg_le_y_old_reg_1 : DFXQD1BWP7T port map(CP => clk, DA => gl_gr_lg_le_y_old(1), DB => sig_logic_y(1), SA => n_0, Q => gl_gr_lg_le_y_old(1));
  gl_gr_lg_le_y_old_reg_0 : DFXQD1BWP7T port map(CP => clk, DA => gl_gr_lg_le_y_old(0), DB => sig_logic_y(0), SA => n_0, Q => gl_gr_lg_le_y_old(0));
  gl_gr_lg_le_y_old_reg_3 : DFXQD1BWP7T port map(CP => clk, DA => gl_gr_lg_le_y_old(3), DB => sig_logic_y(3), SA => n_0, Q => gl_gr_lg_le_y_old(3));
  gl_gr_lg_le_g443 : CKXOR2D1BWP7T port map(A1 => gl_gr_lg_le_x_old(0), A2 => sig_logic_x(0), Z => gl_gr_lg_le_n_7);
  gl_gr_lg_le_g444 : CKXOR2D1BWP7T port map(A1 => gl_gr_lg_le_y_old(2), A2 => sig_logic_y(2), Z => gl_gr_lg_le_n_6);
  gl_gr_lg_le_g445 : CKXOR2D1BWP7T port map(A1 => gl_gr_lg_le_x_old(1), A2 => sig_logic_x(1), Z => gl_gr_lg_le_n_5);
  gl_gr_lg_le_g446 : CKXOR2D1BWP7T port map(A1 => gl_gr_lg_le_y_old(1), A2 => sig_logic_y(1), Z => gl_gr_lg_le_n_4);
  gl_gr_lg_le_g447 : XNR2D1BWP7T port map(A1 => gl_gr_lg_le_y_old(3), A2 => sig_logic_y(3), ZN => gl_gr_lg_le_n_3);
  gl_gr_lg_le_g448 : XNR2D1BWP7T port map(A1 => gl_gr_lg_le_x_old(2), A2 => sig_logic_x(2), ZN => gl_gr_lg_le_n_2);
  gl_gr_lg_le_g449 : XNR2D1BWP7T port map(A1 => gl_gr_lg_le_y_old(0), A2 => sig_logic_y(0), ZN => gl_gr_lg_le_n_1);
  gl_gr_lg_le_g450 : CKXOR2D1BWP7T port map(A1 => gl_gr_lg_le_x_old(3), A2 => sig_logic_x(3), Z => gl_gr_lg_le_n_0);
  gl_gr_lg_lv_count_v_reg_3 : DFQD0BWP7T port map(CP => clk, D => gl_gr_lg_lv_n_15, Q => gl_gr_lg_local_y(3));
  gl_gr_lg_lv_count_v_reg_2 : DFQD0BWP7T port map(CP => clk, D => gl_gr_lg_lv_n_13, Q => gl_gr_lg_local_y(2));
  gl_gr_lg_lv_g403 : OAI31D0BWP7T port map(A1 => gl_gr_lg_lv_n_3, A2 => gl_gr_lg_lv_n_1, A3 => gl_gr_lg_lv_n_6, B => gl_gr_lg_lv_n_14, ZN => gl_gr_lg_lv_n_15);
  gl_gr_lg_lv_g405 : OAI21D0BWP7T port map(A1 => gl_gr_lg_lv_n_10, A2 => gl_gr_lg_lv_n_5, B => gl_gr_lg_local_y(3), ZN => gl_gr_lg_lv_n_14);
  gl_gr_lg_lv_g406 : OAI32D0BWP7T port map(A1 => gl_gr_lg_local_y(2), A2 => gl_gr_lg_lv_n_3, A3 => gl_gr_lg_lv_n_6, B1 => gl_gr_lg_lv_n_1, B2 => gl_gr_lg_lv_n_11, ZN => gl_gr_lg_lv_n_13);
  gl_gr_lg_lv_g407 : OAI22D0BWP7T port map(A1 => gl_gr_lg_lv_n_8, A2 => gl_gr_lg_lv_n_3, B1 => gl_gr_lg_lv_n_6, B2 => gl_gr_lg_local_y(1), ZN => gl_gr_lg_lv_n_12);
  gl_gr_lg_lv_g409 : INVD0BWP7T port map(I => gl_gr_lg_lv_n_10, ZN => gl_gr_lg_lv_n_11);
  gl_gr_lg_lv_g410 : IOA21D1BWP7T port map(A1 => gl_gr_lg_lv_n_5, A2 => gl_gr_lg_lv_n_3, B => gl_gr_lg_lv_n_8, ZN => gl_gr_lg_lv_n_10);
  gl_gr_lg_lv_g412 : AOI21D0BWP7T port map(A1 => gl_gr_lg_lv_n_5, A2 => gl_gr_lg_lv_n_2, B => gl_gr_lg_lv_n_4, ZN => gl_gr_lg_lv_n_8);
  gl_gr_lg_lv_g414 : ND3D0BWP7T port map(A1 => gl_gr_lg_lv_n_5, A2 => gl_gr_lg_lv_sig_edges, A3 => gl_gr_lg_local_y(0), ZN => gl_gr_lg_lv_n_6);
  gl_gr_lg_lv_g415 : AOI31D0BWP7T port map(A1 => gl_gr_lg_local_y(2), A2 => gl_gr_lg_local_y(3), A3 => gl_gr_lg_local_y(1), B => n_0, ZN => gl_gr_lg_lv_n_5);
  gl_gr_lg_lv_g416 : NR2D1BWP7T port map(A1 => gl_gr_lg_lv_sig_edges, A2 => n_0, ZN => gl_gr_lg_lv_n_4);
  gl_gr_lg_lv_fopt422 : INVD0BWP7T port map(I => gl_gr_lg_local_y(2), ZN => gl_gr_lg_lv_n_1);
  gl_gr_lg_lv_count_v_reg_1 : DFD1BWP7T port map(CP => clk, D => gl_gr_lg_lv_n_12, Q => gl_gr_lg_local_y(1), QN => gl_gr_lg_lv_n_3);
  gl_gr_lg_lv_count_v_reg_0 : DFD1BWP7T port map(CP => clk, D => gl_gr_lg_lv_n_19, Q => gl_gr_lg_local_y(0), QN => gl_gr_lg_lv_n_2);
  gl_gr_lg_lv_g2 : AO32D1BWP7T port map(A1 => gl_gr_lg_lv_n_5, A2 => gl_gr_lg_lv_sig_edges, A3 => gl_gr_lg_lv_n_2, B1 => gl_gr_lg_lv_n_4, B2 => gl_gr_lg_local_y(0), Z => gl_gr_lg_lv_n_19);
  gl_gr_lg_lv_l_edge_g12 : NR2XD0BWP7T port map(A1 => gl_gr_lg_lv_l_edge_n_0, A2 => gl_gr_lg_lv_l_edge_reg2, ZN => gl_gr_lg_lv_sig_edges);
  gl_gr_lg_lv_l_edge_reg2_reg : DFQD1BWP7T port map(CP => clk, D => gl_gr_lg_lv_l_edge_reg1, Q => gl_gr_lg_lv_l_edge_reg2);
  gl_gr_lg_lv_l_edge_reg1_reg : DFD1BWP7T port map(CP => clk, D => gl_sig_scale_v, Q => gl_gr_lg_lv_l_edge_reg1, QN => gl_gr_lg_lv_l_edge_n_0);
  ml_ms_ed_reg1_reg : DFQD1BWP7T port map(CP => clk, D => ml_ms_Clk15k_buffered, Q => ml_ms_ed_reg1);
  ml_ms_ed_g247 : NR2XD0BWP7T port map(A1 => ml_ms_ed_n_16, A2 => ml_ms_ed_state(0), ZN => ml_ms_output_edgedet);
  ml_ms_ed_g565 : OAI22D0BWP7T port map(A1 => ml_ms_ed_n_13, A2 => reset, B1 => ml_ms_ed_n_10, B2 => ml_ms_ed_n_6, ZN => ml_ms_ed_n_15);
  ml_ms_ed_g566 : MOAI22D0BWP7T port map(A1 => ml_ms_ed_n_12, A2 => reset, B1 => ml_ms_ed_n_10, B2 => ml_ms_ed_n_0, ZN => ml_ms_ed_n_14);
  ml_ms_ed_g567 : OA31D1BWP7T port map(A1 => ml_ms_ed_reg1, A2 => ml_ms_ed_n_1, A3 => ml_ms_ed_state(0), B => ml_ms_ed_n_12, Z => ml_ms_ed_n_13);
  ml_ms_ed_g568 : OA21D0BWP7T port map(A1 => ml_ms_ed_n_16, A2 => ml_ms_ed_state(0), B => ml_ms_ed_n_35, Z => ml_ms_ed_n_12);
  ml_ms_ed_g570 : ND3D0BWP7T port map(A1 => ml_ms_ed_n_9, A2 => ml_ms_ed_n_7, A3 => ml_ms_ed_n_5, ZN => ml_ms_ed_n_10);
  ml_ms_ed_g571 : OAI31D0BWP7T port map(A1 => ml_ms_count_debounce(6), A2 => ml_ms_count_debounce(5), A3 => ml_ms_ed_n_4, B => ml_ms_count_debounce(7), ZN => ml_ms_ed_n_9);
  ml_ms_ed_g572 : IND4D0BWP7T port map(A1 => ml_ms_ed_n_5, B1 => ml_ms_count_debounce(5), B2 => ml_ms_count_debounce(6), B3 => ml_ms_ed_n_3, ZN => ml_ms_ed_n_8);
  ml_ms_ed_g573 : NR4D0BWP7T port map(A1 => ml_ms_ed_n_2, A2 => ml_ms_count_debounce(12), A3 => ml_ms_count_debounce(9), A4 => ml_ms_count_debounce(10), ZN => ml_ms_ed_n_7);
  ml_ms_ed_g574 : INVD1BWP7T port map(I => ml_ms_ed_n_0, ZN => ml_ms_ed_n_6);
  ml_ms_ed_g576 : AN3D0BWP7T port map(A1 => ml_ms_count_debounce(2), A2 => ml_ms_count_debounce(4), A3 => ml_ms_count_debounce(1), Z => ml_ms_ed_n_4);
  ml_ms_ed_g577 : ND3D0BWP7T port map(A1 => ml_ms_count_debounce(7), A2 => ml_ms_count_debounce(4), A3 => ml_ms_count_debounce(3), ZN => ml_ms_ed_n_5);
  ml_ms_ed_g578 : OR2D1BWP7T port map(A1 => ml_ms_count_debounce(1), A2 => ml_ms_count_debounce(2), Z => ml_ms_ed_n_3);
  ml_ms_ed_g579 : OR2D1BWP7T port map(A1 => ml_ms_count_debounce(11), A2 => ml_ms_count_debounce(8), Z => ml_ms_ed_n_2);
  ml_ms_ed_g2 : INR3D0BWP7T port map(A1 => ml_ms_ed_state(0), B1 => ml_ms_ed_state(1), B2 => reset, ZN => ml_ms_ed_n_0);
  ml_ms_ed_g586 : ND3D0BWP7T port map(A1 => ml_ms_ed_n_8, A2 => ml_ms_ed_n_7, A3 => ml_ms_ed_state(1), ZN => ml_ms_ed_n_35);
  ml_ms_ed_state_reg_0 : DFD1BWP7T port map(CP => clk, D => ml_ms_ed_n_15, Q => ml_ms_ed_state(0), QN => ml_ms_count_debounce_reset);
  ml_ms_ed_state_reg_1 : DFD1BWP7T port map(CP => clk, D => ml_ms_ed_n_14, Q => ml_ms_ed_state(1), QN => ml_ms_ed_n_16);
  ml_ms_ed_reg2_reg : DFD1BWP7T port map(CP => clk, D => ml_ms_ed_reg1, Q => ml_ms_ed_reg2, QN => ml_ms_ed_n_1);
  ml_ms_cntD_g71 : INVD1BWP7T port map(I => ml_ms_count_debounce_reset, ZN => ml_ms_cntD_n_23);
  ml_ms_cntD_count_reg_12 : DFKCNQD1BWP7T port map(CP => clk, CN => ml_ms_cntD_n_23, D => ml_ms_cntD_n_22, Q => ml_ms_count_debounce(12));
  ml_ms_cntD_count_reg_11 : DFKCNQD1BWP7T port map(CP => clk, CN => ml_ms_cntD_n_23, D => ml_ms_cntD_n_21, Q => ml_ms_count_debounce(11));
  ml_ms_cntD_g225 : MOAI22D0BWP7T port map(A1 => ml_ms_cntD_n_20, A2 => ml_ms_count_debounce(12), B1 => ml_ms_cntD_n_20, B2 => ml_ms_count_debounce(12), ZN => ml_ms_cntD_n_22);
  ml_ms_cntD_count_reg_10 : DFKCNQD1BWP7T port map(CP => clk, CN => ml_ms_cntD_n_23, D => ml_ms_cntD_n_19, Q => ml_ms_count_debounce(10));
  ml_ms_cntD_g227 : MOAI22D0BWP7T port map(A1 => ml_ms_cntD_n_18, A2 => ml_ms_count_debounce(11), B1 => ml_ms_cntD_n_18, B2 => ml_ms_count_debounce(11), ZN => ml_ms_cntD_n_21);
  ml_ms_cntD_g228 : IND2D1BWP7T port map(A1 => ml_ms_cntD_n_18, B1 => ml_ms_count_debounce(11), ZN => ml_ms_cntD_n_20);
  ml_ms_cntD_count_reg_9 : DFKCNQD1BWP7T port map(CP => clk, CN => ml_ms_cntD_n_23, D => ml_ms_cntD_n_17, Q => ml_ms_count_debounce(9));
  ml_ms_cntD_g230 : MOAI22D0BWP7T port map(A1 => ml_ms_cntD_n_16, A2 => ml_ms_count_debounce(10), B1 => ml_ms_cntD_n_16, B2 => ml_ms_count_debounce(10), ZN => ml_ms_cntD_n_19);
  ml_ms_cntD_g231 : IND2D1BWP7T port map(A1 => ml_ms_cntD_n_16, B1 => ml_ms_count_debounce(10), ZN => ml_ms_cntD_n_18);
  ml_ms_cntD_count_reg_8 : DFKCNQD1BWP7T port map(CP => clk, CN => ml_ms_cntD_n_23, D => ml_ms_cntD_n_15, Q => ml_ms_count_debounce(8));
  ml_ms_cntD_g233 : MOAI22D0BWP7T port map(A1 => ml_ms_cntD_n_14, A2 => ml_ms_count_debounce(9), B1 => ml_ms_cntD_n_14, B2 => ml_ms_count_debounce(9), ZN => ml_ms_cntD_n_17);
  ml_ms_cntD_g234 : IND2D1BWP7T port map(A1 => ml_ms_cntD_n_14, B1 => ml_ms_count_debounce(9), ZN => ml_ms_cntD_n_16);
  ml_ms_cntD_count_reg_7 : DFKCNQD1BWP7T port map(CP => clk, CN => ml_ms_cntD_n_23, D => ml_ms_cntD_n_13, Q => ml_ms_count_debounce(7));
  ml_ms_cntD_g236 : MOAI22D0BWP7T port map(A1 => ml_ms_cntD_n_12, A2 => ml_ms_count_debounce(8), B1 => ml_ms_cntD_n_12, B2 => ml_ms_count_debounce(8), ZN => ml_ms_cntD_n_15);
  ml_ms_cntD_g237 : IND2D1BWP7T port map(A1 => ml_ms_cntD_n_12, B1 => ml_ms_count_debounce(8), ZN => ml_ms_cntD_n_14);
  ml_ms_cntD_count_reg_6 : DFKCNQD1BWP7T port map(CP => clk, CN => ml_ms_cntD_n_23, D => ml_ms_cntD_n_11, Q => ml_ms_count_debounce(6));
  ml_ms_cntD_g239 : MOAI22D0BWP7T port map(A1 => ml_ms_cntD_n_10, A2 => ml_ms_count_debounce(7), B1 => ml_ms_cntD_n_10, B2 => ml_ms_count_debounce(7), ZN => ml_ms_cntD_n_13);
  ml_ms_cntD_g240 : IND2D1BWP7T port map(A1 => ml_ms_cntD_n_10, B1 => ml_ms_count_debounce(7), ZN => ml_ms_cntD_n_12);
  ml_ms_cntD_count_reg_5 : DFKCNQD1BWP7T port map(CP => clk, CN => ml_ms_cntD_n_23, D => ml_ms_cntD_n_9, Q => ml_ms_count_debounce(5));
  ml_ms_cntD_g242 : MOAI22D0BWP7T port map(A1 => ml_ms_cntD_n_8, A2 => ml_ms_count_debounce(6), B1 => ml_ms_cntD_n_8, B2 => ml_ms_count_debounce(6), ZN => ml_ms_cntD_n_11);
  ml_ms_cntD_g243 : IND2D1BWP7T port map(A1 => ml_ms_cntD_n_8, B1 => ml_ms_count_debounce(6), ZN => ml_ms_cntD_n_10);
  ml_ms_cntD_count_reg_4 : DFKCNQD1BWP7T port map(CP => clk, CN => ml_ms_cntD_n_23, D => ml_ms_cntD_n_7, Q => ml_ms_count_debounce(4));
  ml_ms_cntD_g245 : MOAI22D0BWP7T port map(A1 => ml_ms_cntD_n_6, A2 => ml_ms_count_debounce(5), B1 => ml_ms_cntD_n_6, B2 => ml_ms_count_debounce(5), ZN => ml_ms_cntD_n_9);
  ml_ms_cntD_g246 : IND2D1BWP7T port map(A1 => ml_ms_cntD_n_6, B1 => ml_ms_count_debounce(5), ZN => ml_ms_cntD_n_8);
  ml_ms_cntD_count_reg_3 : DFKCNQD1BWP7T port map(CP => clk, CN => ml_ms_cntD_n_23, D => ml_ms_cntD_n_5, Q => ml_ms_count_debounce(3));
  ml_ms_cntD_g248 : MOAI22D0BWP7T port map(A1 => ml_ms_cntD_n_4, A2 => ml_ms_count_debounce(4), B1 => ml_ms_cntD_n_4, B2 => ml_ms_count_debounce(4), ZN => ml_ms_cntD_n_7);
  ml_ms_cntD_g249 : IND2D1BWP7T port map(A1 => ml_ms_cntD_n_4, B1 => ml_ms_count_debounce(4), ZN => ml_ms_cntD_n_6);
  ml_ms_cntD_count_reg_2 : DFKCNQD1BWP7T port map(CP => clk, CN => ml_ms_cntD_n_23, D => ml_ms_cntD_n_3, Q => ml_ms_count_debounce(2));
  ml_ms_cntD_g251 : MOAI22D0BWP7T port map(A1 => ml_ms_cntD_n_2, A2 => ml_ms_count_debounce(3), B1 => ml_ms_cntD_n_2, B2 => ml_ms_count_debounce(3), ZN => ml_ms_cntD_n_5);
  ml_ms_cntD_g252 : IND2D1BWP7T port map(A1 => ml_ms_cntD_n_2, B1 => ml_ms_count_debounce(3), ZN => ml_ms_cntD_n_4);
  ml_ms_cntD_count_reg_1 : DFKCNQD1BWP7T port map(CP => clk, CN => ml_ms_cntD_n_23, D => ml_ms_cntD_n_1, Q => ml_ms_count_debounce(1));
  ml_ms_cntD_g254 : MOAI22D0BWP7T port map(A1 => ml_ms_cntD_n_0, A2 => ml_ms_count_debounce(2), B1 => ml_ms_cntD_n_0, B2 => ml_ms_count_debounce(2), ZN => ml_ms_cntD_n_3);
  ml_ms_cntD_g255 : IND2D1BWP7T port map(A1 => ml_ms_cntD_n_0, B1 => ml_ms_count_debounce(2), ZN => ml_ms_cntD_n_2);
  ml_ms_cntD_count_reg_0 : DFKCND1BWP7T port map(CP => clk, CN => ml_ms_cntD_count(0), D => ml_ms_cntD_n_23, Q => UNCONNECTED2, QN => ml_ms_cntD_count(0));
  ml_ms_cntD_g257 : MOAI22D0BWP7T port map(A1 => ml_ms_cntD_count(0), A2 => ml_ms_count_debounce(1), B1 => ml_ms_cntD_count(0), B2 => ml_ms_count_debounce(1), ZN => ml_ms_cntD_n_1);
  ml_ms_cntD_g258 : IND2D1BWP7T port map(A1 => ml_ms_cntD_count(0), B1 => ml_ms_count_debounce(1), ZN => ml_ms_cntD_n_0);
  gl_gr_lg_lh_count_h_reg_3 : DFQD0BWP7T port map(CP => clk, D => gl_gr_lg_lh_n_15, Q => gl_gr_lg_local_x(3));
  gl_gr_lg_lh_g403 : OAI31D0BWP7T port map(A1 => gl_gr_lg_lh_n_3, A2 => gl_gr_lg_lh_n_1, A3 => gl_gr_lg_lh_n_6, B => gl_gr_lg_lh_n_14, ZN => gl_gr_lg_lh_n_15);
  gl_gr_lg_lh_g405 : OAI21D0BWP7T port map(A1 => gl_gr_lg_lh_n_10, A2 => gl_gr_lg_lh_n_5, B => gl_gr_lg_local_x(3), ZN => gl_gr_lg_lh_n_14);
  gl_gr_lg_lh_g406 : OAI32D0BWP7T port map(A1 => gl_gr_lg_local_x(2), A2 => gl_gr_lg_lh_n_3, A3 => gl_gr_lg_lh_n_6, B1 => gl_gr_lg_lh_n_1, B2 => gl_gr_lg_lh_n_11, ZN => gl_gr_lg_lh_n_13);
  gl_gr_lg_lh_g407 : OAI22D0BWP7T port map(A1 => gl_gr_lg_lh_n_8, A2 => gl_gr_lg_lh_n_3, B1 => gl_gr_lg_lh_n_6, B2 => gl_gr_lg_local_x(1), ZN => gl_gr_lg_lh_n_12);
  gl_gr_lg_lh_g409 : INVD0BWP7T port map(I => gl_gr_lg_lh_n_10, ZN => gl_gr_lg_lh_n_11);
  gl_gr_lg_lh_g410 : IOA21D1BWP7T port map(A1 => gl_gr_lg_lh_n_5, A2 => gl_gr_lg_lh_n_3, B => gl_gr_lg_lh_n_8, ZN => gl_gr_lg_lh_n_10);
  gl_gr_lg_lh_g412 : AOI21D0BWP7T port map(A1 => gl_gr_lg_lh_n_5, A2 => gl_gr_lg_lh_n_2, B => gl_gr_lg_lh_n_4, ZN => gl_gr_lg_lh_n_8);
  gl_gr_lg_lh_g414 : ND3D0BWP7T port map(A1 => gl_gr_lg_lh_n_5, A2 => gl_gr_lg_lh_sig_edges, A3 => gl_gr_lg_local_x(0), ZN => gl_gr_lg_lh_n_6);
  gl_gr_lg_lh_g415 : AOI31D0BWP7T port map(A1 => gl_gr_lg_local_x(2), A2 => gl_gr_lg_local_x(3), A3 => gl_gr_lg_local_x(1), B => n_0, ZN => gl_gr_lg_lh_n_5);
  gl_gr_lg_lh_g416 : NR2D1BWP7T port map(A1 => gl_gr_lg_lh_sig_edges, A2 => n_0, ZN => gl_gr_lg_lh_n_4);
  gl_gr_lg_lh_count_h_reg_1 : DFD1BWP7T port map(CP => clk, D => gl_gr_lg_lh_n_12, Q => gl_gr_lg_local_x(1), QN => gl_gr_lg_lh_n_3);
  gl_gr_lg_lh_count_h_reg_0 : DFD1BWP7T port map(CP => clk, D => gl_gr_lg_lh_n_19, Q => gl_gr_lg_local_x(0), QN => gl_gr_lg_lh_n_2);
  gl_gr_lg_lh_count_h_reg_2 : DFD1BWP7T port map(CP => clk, D => gl_gr_lg_lh_n_13, Q => gl_gr_lg_local_x(2), QN => gl_gr_lg_lh_n_1);
  gl_gr_lg_lh_g2 : AO32D1BWP7T port map(A1 => gl_gr_lg_lh_n_5, A2 => gl_gr_lg_lh_sig_edges, A3 => gl_gr_lg_lh_n_2, B1 => gl_gr_lg_lh_n_4, B2 => gl_gr_lg_local_x(0), Z => gl_gr_lg_lh_n_19);
  gl_gr_lg_lh_l_edge_g12 : NR2XD0BWP7T port map(A1 => gl_gr_lg_lh_l_edge_n_0, A2 => gl_gr_lg_lh_l_edge_reg2, ZN => gl_gr_lg_lh_sig_edges);
  gl_gr_lg_lh_l_edge_reg2_reg : DFQD1BWP7T port map(CP => clk, D => gl_gr_lg_lh_l_edge_reg1, Q => gl_gr_lg_lh_l_edge_reg2);
  gl_gr_lg_lh_l_edge_reg1_reg : DFD1BWP7T port map(CP => clk, D => gl_sig_scale_h, Q => gl_gr_lg_lh_l_edge_reg1, QN => gl_gr_lg_lh_l_edge_n_0);

end synthesised;
