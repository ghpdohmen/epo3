
library ieee;
use ieee.std_logic_1164.all;
--library tcb018gbwp7t;
--use tcb018gbwp7t.all;

architecture routed of pixel is

  component BUFFD1P5BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL01BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL02BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component BUFFD3BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKBD0BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component BUFFD2BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKBD2BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL015BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component BUFFD0BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL0BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKBD3BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component BUFFD5BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL1BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component DEL2BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component INVD1BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component CKND2BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component CKBD10BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component INVD2BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component HA1D0BWP7T
    port(A, B : in std_logic; CO, S : out std_logic);
  end component;

  component AO21D0BWP7T
    port(A1, A2, B : in std_logic; Z : out std_logic);
  end component;

  component NR2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component MOAI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component CKXOR2D0BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component AOI21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component MAOI222D0BWP7T
    port(A, B, C : in std_logic; ZN : out std_logic);
  end component;

  component IND2D0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component INR2D0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component ND2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component CKND1BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component ND2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component AOI222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; ZN : out std_logic);
  end component;

  component NR3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component IND3D1BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component INR3D0BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component ND4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component DFKCNQD1BWP7T
    port(CN, CP, D : in std_logic; Q : out std_logic);
  end component;

  component INR4D0BWP7T
    port(A1, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component DFD1BWP7T
    port(CP, D : in std_logic; Q, QN : out std_logic);
  end component;

  component LNQD1BWP7T
    port(D, EN : in std_logic; Q : out std_logic);
  end component;

  component AN3D0BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component NR4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component OAI211D1BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component NR2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component AOI211XD0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component AN4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component XNR2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component CKXOR2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component CKAN2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component OR2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component IND2D1BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component CKND2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component INVD0BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component MAOI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AO32D1BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component IINR4D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI32D1BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AOI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component CKND2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component INR2XD0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component OA21D0BWP7T
    port(A1, A2, B : in std_logic; Z : out std_logic);
  end component;

  component NR2XD0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component AN2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component INR2D1BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component LHQD1BWP7T
    port(D, E : in std_logic; Q : out std_logic);
  end component;

  component NR2XD1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component INR2D2BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component AN2D2BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component AN4D1BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component FA1D0BWP7T
    port(A, B, CI : in std_logic; CO, S : out std_logic);
  end component;

  component DFQD1BWP7T
    port(CP, D : in std_logic; Q : out std_logic);
  end component;

  component OAI31D0BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component AOI221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; ZN : out std_logic);
  end component;

  component AO221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; Z : out std_logic);
  end component;

  component OAI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AOI31D0BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component OAI222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; ZN : out std_logic);
  end component;

  component AO222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; Z : out std_logic);
  end component;

  component AOI33D1BWP7T
    port(A1, A2, A3, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component AO211D0BWP7T
    port(A1, A2, B, C : in std_logic; Z : out std_logic);
  end component;

  component IOA21D1BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component AN2D0BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component AO22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component NR2D1P5BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component OA211D0BWP7T
    port(A1, A2, B, C : in std_logic; Z : out std_logic);
  end component;

  component AN3D1BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component NR3D1BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component ND3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component OR3D1BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component OR2D2BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component DFD0BWP7T
    port(CP, D : in std_logic; Q, QN : out std_logic);
  end component;

  component EDFQD1BWP7T
    port(CP, D, E : in std_logic; Q : out std_logic);
  end component;

  component EDFQD0BWP7T
    port(CP, D, E : in std_logic; Q : out std_logic);
  end component;

  component AOI21D2BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component DFQD0BWP7T
    port(CP, D : in std_logic; Q : out std_logic);
  end component;

  component OAI32D0BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component IAO21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component OA31D1BWP7T
    port(A1, A2, A3, B : in std_logic; Z : out std_logic);
  end component;

  component OA22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component IND4D0BWP7T
    port(A1, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component OAI31D1BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component OR4D1BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component EDFKCNQD1BWP7T
    port(CN, CP, D, E : in std_logic; Q : out std_logic);
  end component;

  component CKXOR2D2BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component DFXQD1BWP7T
    port(CP, DA, DB, SA : in std_logic; Q : out std_logic);
  end component;

  component EDFKCND1BWP7T
    port(CN, CP, D, E : in std_logic; Q, QN : out std_logic);
  end component;

  component DFKCND1BWP7T
    port(CN, CP, D : in std_logic; Q, QN : out std_logic);
  end component;

  component ND2D5BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component MUX2D1BWP7T
    port(I0, I1, S : in std_logic; Z : out std_logic);
  end component;

  component OA32D1BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component MUX2ND0BWP7T
    port(I0, I1, S : in std_logic; ZN : out std_logic);
  end component;

  component IIND4D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AOI32D1BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OA222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; Z : out std_logic);
  end component;

  signal FE_PHN672_gl_ram_n_470, FE_PHN671_gl_ram_n_435, FE_PHN670_gl_ram_ram_35_0, FE_PHN669_gl_ram_ram_27_2, FE_PHN668_gl_ram_ram_1_2 : std_logic;
  signal FE_PHN667_gl_ram_ram_33_0, FE_PHN666_ml_ms_count_debounce_12, FE_PHN665_gl_ram_ram_21_0, FE_PHN664_gl_ram_ram_58_1, FE_PHN663_ml_ms_count_debounce_12 : std_logic;
  signal FE_PHN662_gl_ram_ram_37_2, FE_PHN661_gl_ram_ram_75_0, FE_PHN660_gl_ram_ram_59_2, FE_PHN659_gl_ram_ram_18_0, FE_PHN658_gl_ram_ram_43_1 : std_logic;
  signal FE_PHN657_gl_ram_n_445, FE_PHN656_ml_ms_ed_n_8, FE_PHN655_ml_ms_count_debounce_7, FE_PHN654_gl_ram_ram_17_1, FE_PHN653_ml_ms_count_debounce_12 : std_logic;
  signal FE_PHN652_gl_ram_ram_11_2, FE_PHN651_gl_ram_ram_16_2, FE_PHN650_gl_ram_ram_97_1, FE_PHN649_gl_ram_ram_34_1, FE_PHN648_gl_ram_ram_9_2 : std_logic;
  signal FE_PHN647_gl_ram_ram_8_1, FE_PHN646_gl_ram_ram_8_2, FE_PHN645_gl_ram_ram_51_2, FE_PHN644_gl_ram_ram_12_2, FE_PHN643_gl_ram_ram_88_0 : std_logic;
  signal FE_PHN642_gl_ram_ram_12_1, FE_PHN641_ml_ms_sr_new_new_data_4, FE_PHN640_gl_ram_ram_91_1, FE_PHN639_gl_ram_ram_27_0, FE_PHN638_gl_ram_ram_5_1 : std_logic;
  signal FE_PHN637_gl_ram_ram_48_1, FE_PHN636_ml_ms_ed_reg2, FE_PHN635_gl_ram_ram_27_2, FE_PHN634_gl_ram_ram_50_2, FE_PHN633_gl_ram_ram_50_1 : std_logic;
  signal FE_PHN632_gl_ram_ram_57_1, FE_PHN631_gl_ram_ram_33_2, FE_PHN630_gl_ram_ram_25_0, FE_PHN629_gl_ram_ram_29_1, FE_PHN628_gl_ram_n_437 : std_logic;
  signal FE_PHN627_gl_ram_n_523, FE_PHN626_gl_ram_ram_41_0, FE_PHN625_gl_ram_ram_4_0, FE_PHN624_gl_ram_ram_89_0, FE_PHN623_ml_ms_sr_new_new_data_0 : std_logic;
  signal FE_PHN622_ml_ms_ed_n_8, FE_PHN621_ml_ms_ed_n_2, FE_PHN620_ml_ms_n_23, FE_PHN619_ml_ms_n_24, FE_PHN618_ml_ms_n_22 : std_logic;
  signal FE_PHN617_ml_ms_count_debounce_10, FE_PHN616_ml_ms_count_debounce_6, FE_PHN615_ml_ms_count_debounce_12, FE_PHN614_ml_ms_ed_state_0, FE_PHN613_ml_ms_sr_new_new_data_0 : std_logic;
  signal FE_PHN612_ml_ms_count_debounce_7, FE_PHN611_gl_ram_ram_19_1, FE_PHN610_ml_ms_ed_state_1, FE_PHN609_gl_ram_ram_17_1, FE_PHN608_gl_ram_ram_97_1 : std_logic;
  signal FE_PHN607_gl_ram_ram_12_2, FE_PHN606_gl_ram_ram_58_1, FE_PHN605_gl_ram_ram_24_2, FE_PHN604_gl_ram_ram_73_2, FE_PHN603_gl_ram_ram_4_0 : std_logic;
  signal FE_PHN602_gl_ram_ram_88_0, FE_PHN601_gl_ram_ram_21_0, FE_PHN600_gl_ram_ram_32_1, FE_PHN599_gl_ram_ram_18_0, FE_PHN598_gl_ram_ram_16_2 : std_logic;
  signal FE_PHN597_gl_ram_ram_2_2, FE_PHN596_gl_ram_ram_27_0, FE_PHN595_gl_ram_ram_12_1, FE_PHN594_gl_ram_ram_89_0, FE_PHN593_gl_ram_ram_37_2 : std_logic;
  signal FE_PHN592_gl_ram_ram_35_2, FE_PHN591_gl_ram_ram_56_2, FE_PHN590_gl_ram_ram_56_1, FE_PHN589_gl_ram_ram_50_2, FE_PHN588_gl_ram_ram_50_1 : std_logic;
  signal FE_PHN587_gl_ram_ram_29_1, FE_PHN586_gl_ram_ram_51_2, FE_PHN585_gl_ram_ram_33_0, FE_PHN584_gl_ram_ram_48_1, FE_PHN583_gl_ram_ram_35_0 : std_logic;
  signal FE_PHN582_gl_ram_ram_41_0, FE_PHN581_gl_ram_ram_57_1, FE_PHN580_gl_ram_ram_75_0, FE_PHN579_gl_ram_n_489, FE_PHN578_gl_ram_ram_8_2 : std_logic;
  signal FE_PHN577_gl_ram_ram_25_0, FE_PHN576_gl_ram_ram_33_2, FE_PHN575_gl_ram_ram_8_0, FE_PHN574_gl_ram_ram_91_1, FE_PHN573_gl_ram_ram_11_2 : std_logic;
  signal FE_PHN572_gl_ram_ram_8_1, FE_PHN571_gl_ram_ram_34_1, FE_PHN570_gl_ram_ram_82_0, FE_PHN569_gl_ram_ram_2_0, FE_PHN568_gl_ram_ram_11_1 : std_logic;
  signal FE_PHN567_gl_ram_ram_3_2, FE_PHN566_ml_ms_muxReg, FE_PHN565_gl_ram_ram_9_0, FE_PHN564_gl_ram_ram_43_2, FE_PHN563_gl_ram_ram_24_0 : std_logic;
  signal FE_PHN562_gl_ram_ram_3_0, FE_PHN561_gl_ram_ram_1_0, FE_PHN560_gl_ram_ram_0_1, FE_PHN559_gl_ram_ram_43_0, FE_PHN558_gl_ram_ram_19_0 : std_logic;
  signal FE_PHN557_gl_ram_ram_24_1, FE_PHN556_gl_ram_ram_32_0, FE_PHN555_gl_ram_ram_27_1, FE_PHN554_gl_ram_ram_40_0, FE_PHN553_gl_ram_ram_0_0 : std_logic;
  signal FE_PHN552_ml_ms_sr_new_new_data_6, FE_PHN551_ml_ms_ed_n_8, FE_PHN550_ml_ms_n_34, FE_PHN549_ml_ms_n_32, FE_PHN548_ml_ms_n_30 : std_logic;
  signal FE_PHN547_ml_ms_ed_n_5, FE_PHN546_ml_ms_n_58, FE_PHN545_ml_ms_n_21, FE_PHN544_ml_ms_n_60, FE_PHN543_gl_vgd_horizontal_counter_6 : std_logic;
  signal FE_PHN542_ml_ms_data_sr_11bit_3, FE_PHN541_gl_ram_ram_8_2, FE_PHN540_gl_ram_ram_25_0, FE_PHN539_gl_ram_ram_57_1, FE_PHN538_gl_ram_ram_19_0 : std_logic;
  signal FE_PHN537_gl_ram_ram_50_2, FE_PHN536_gl_ram_ram_41_0, FE_PHN535_gl_ram_ram_12_2, FE_PHN534_gl_ram_ram_8_1, FE_PHN533_gl_ram_ram_48_2 : std_logic;
  signal FE_PHN532_gl_ram_ram_11_0, FE_PHN531_gl_ram_ram_89_0, FE_PHN530_gl_ram_ram_27_0, FE_PHN529_gl_vgd_horizontal_counter_7, FE_PHN528_gl_ram_ram_9_2 : std_logic;
  signal FE_PHN527_gl_ram_ram_40_1, FE_PHN526_ml_ms_muxFSM, FE_PHN525_gl_ram_ram_43_1, FE_PHN524_gl_vgd_horizontal_counter_8, FE_PHN523_gl_ram_ram_0_2 : std_logic;
  signal FE_PHN522_gl_ram_ram_21_0, FE_PHN521_gl_ram_ram_24_2, FE_PHN520_gl_ram_ram_58_1, FE_PHN519_gl_ram_ram_1_2, FE_PHN518_gl_ram_ram_27_2 : std_logic;
  signal FE_PHN517_gl_ram_ram_2_2, FE_PHN516_ml_ms_sr_new_new_data_5, FE_PHN515_ml_ms_sfsm_state_0, FE_PHN514_gl_ram_ram_88_0, FE_PHN513_ml_ms_count_debounce_6 : std_logic;
  signal FE_PHN512_gl_ram_ram_43_2, FE_PHN511_gl_ram_ram_17_1, FE_PHN510_gl_ram_ram_11_2, FE_PHN509_gl_ram_ram_37_2, FE_PHN508_gl_ram_ram_11_1 : std_logic;
  signal FE_PHN507_gl_ram_ram_4_0, FE_PHN506_gl_ram_ram_0_1, FE_PHN505_gl_ram_ram_2_0, FE_PHN504_gl_ram_ram_12_1, FE_PHN503_gl_ram_ram_3_2 : std_logic;
  signal FE_PHN502_gl_ram_ram_51_2, FE_PHN501_gl_ram_ram_56_1, FE_PHN500_gl_ram_ram_56_2, FE_PHN499_gl_ram_ram_8_0, FE_PHN498_gl_ram_ram_75_0 : std_logic;
  signal FE_PHN497_gl_ram_ram_32_1, FE_PHN496_gl_ram_ram_24_0, FE_PHN495_gl_ram_ram_29_1, FE_PHN494_gl_ram_ram_43_0, FE_PHN493_gl_ram_ram_35_0 : std_logic;
  signal FE_PHN492_gl_ram_ram_5_1, FE_PHN491_gl_ram_ram_9_0, FE_PHN490_gl_ram_ram_48_1, FE_PHN489_gl_ram_ram_1_0, FE_PHN488_gl_ram_ram_33_0 : std_logic;
  signal FE_PHN487_gl_ram_ram_3_0, FE_PHN486_gl_ram_ram_24_1, FE_PHN485_gl_ram_ram_59_2, FE_PHN484_gl_ram_ram_40_0, FE_PHN483_gl_ram_ram_32_0 : std_logic;
  signal FE_PHN482_gl_ram_ram_33_2, FE_PHN481_gl_ram_ram_0_0, FE_PHN480_gl_ram_ram_97_1, FE_PHN479_gl_ram_ram_91_1, FE_PHN478_gl_ram_ram_27_1 : std_logic;
  signal FE_PHN477_gl_ram_ram_35_2, FE_PHN476_gl_ram_ram_19_1, FE_PHN475_gl_ram_ram_34_1, FE_PHN474_gl_ram_ram_50_1, FE_PHN473_ml_ms_count_debounce_7 : std_logic;
  signal FE_PHN472_gl_ram_ram_73_2, FE_PHN471_gl_ram_n_396, FE_PHN470_ml_ms_ed_n_2, FE_PHN469_gl_ram_n_400, FE_PHN468_ml_ms_sr_new_new_data_6 : std_logic;
  signal FE_PHN467_ml_ms_mfsm_n_21, FE_PHN466_ml_ms_sr_new_new_data_7, FE_PHN465_gl_gr_lg_local_y_0, FE_PHN464_sig_logic_y_0, FE_PHN463_ml_ms_count_debounce_10 : std_logic;
  signal FE_PHN462_gl_ram_ram_82_0, FE_PHN461_ml_il_color1_n_15, FE_PHN460_ml_ms_n_31, FE_PHN459_ml_ms_n_24, FE_PHN458_ml_ms_n_60 : std_logic;
  signal FE_PHN457_ml_ms_n_58, FE_PHN456_ml_ms_mfsm_n_52, FE_PHN455_gl_gr_lg_lv_n_15, FE_PHN454_ml_ms_mfsm_n_0, FE_PHN453_gl_vgd_horizontal_counter_6 : std_logic;
  signal FE_PHN452_ml_ms_count25M_8, FE_PHN451_gl_ram_ram_82_0, FE_PHN450_gl_ram_ram_20_2, FE_PHN449_gl_ram_ram_46_2, FE_PHN448_ml_ms_tb_n_0 : std_logic;
  signal FE_PHN447_gl_ram_ram_37_0, FE_PHN446_ml_ms_mux_select, FE_PHN445_gl_gr_lg_lcountdown_n_2, FE_PHN444_gl_ram_ram_80_0, FE_PHN443_gl_gr_lg_lcountdown_n_4 : std_logic;
  signal FE_PHN442_gl_ram_ram_5_0, FE_PHN441_ml_ms_n_2, FE_PHN440_gl_ram_ram_86_1, FE_PHN439_gl_ram_ram_61_1, FE_PHN438_gl_ram_ram_10_0 : std_logic;
  signal FE_PHN437_ml_il_color1_n_15, FE_PHN436_sig_logic_y_0, FE_PHN435_gl_gr_lg_lcountdown_n_15, FE_PHN434_ml_ms_count_debounce_6, FE_PHN433_ml_ms_count_debounce_10 : std_logic;
  signal FE_PHN432_ml_ms_data_sr_11bit_3, FE_PHN431_gl_ram_ram_60_0, FE_PHN430_gl_ram_ram_60_2, FE_PHN429_gl_ram_ram_60_1, FE_PHN428_gl_ram_ram_36_2 : std_logic;
  signal FE_PHN427_gl_ram_ram_33_1, FE_PHN426_gl_ram_ram_96_2, FE_PHN425_gl_ram_n_495, FE_PHN424_gl_ram_ram_31_2, FE_PHN423_gl_ram_ram_25_1 : std_logic;
  signal FE_PHN422_gl_ram_ram_20_1, FE_PHN421_gl_ram_ram_65_2, FE_PHN420_gl_ram_ram_97_0, FE_PHN419_gl_ram_ram_96_1, FE_PHN418_gl_ram_ram_83_0 : std_logic;
  signal FE_PHN417_gl_ram_ram_73_0, FE_PHN416_gl_ram_ram_66_0, FE_PHN415_gl_ram_n_496, FE_PHN414_gl_ram_ram_67_0, FE_PHN413_gl_ram_n_394 : std_logic;
  signal FE_PHN412_gl_ram_ram_73_1, FE_PHN411_gl_ram_ram_41_2, FE_PHN410_ml_ms_cnt_count_0, FE_PHN409_gl_ram_ram_98_2, FE_PHN408_gl_ram_ram_82_1 : std_logic;
  signal FE_PHN407_gl_gr_lg_lv_n_3, FE_PHN406_ml_il_color1_state_hs_1, FE_PHN405_gl_gr_lg_lcountdown_n_13, FE_PHN404_gl_gr_lg_lcountdown_n_17, FE_PHN403_gl_gr_lg_lcountdown_n_19 : std_logic;
  signal FE_PHN402_gl_gr_lg_lcountdown_n_8, FE_PHN401_gl_gr_lg_lcountdown_n_20, FE_PHN400_gl_gr_lg_lcountdown_n_11, FE_PHN399_gl_gr_lg_lcountdown_n_21, FE_PHN398_gl_gr_lg_lcountdown_n_0 : std_logic;
  signal FE_PHN397_ml_ms_cntD_n_19, FE_PHN396_gl_gr_lg_lcountdown_sig_edge_fall, FE_PHN395_ml_il_x1_n_9, FE_PHN394_ml_ms_mfsm_n_44, FE_PHN393_ml_ms_cnt_n_5 : std_logic;
  signal FE_PHN392_gl_ram_n_145, FE_PHN391_ml_ms_tb_n_5, FE_PHN390_ml_ms_cnt_n_9, FE_PHN389_gl_ram_n_563, FE_PHN388_ml_ms_tb_n_6 : std_logic;
  signal FE_PHN387_ml_ms_mfsm_n_38, FE_PHN386_ml_ms_cnt_n_7, FE_PHN385_ml_il_color1_n_14, FE_PHN384_ml_il_y1_n_9, FE_PHN383_ml_ms_cnt_n_3 : std_logic;
  signal FE_PHN382_gl_ram_n_564, FE_PHN381_gl_ram_n_567, FE_PHN380_gl_gr_lg_lv_n_12, FE_PHN379_ml_ms_n_54, FE_PHN378_ml_il_color1_n_13 : std_logic;
  signal FE_PHN377_gl_ram_n_247, FE_PHN376_gl_ram_n_308, FE_PHN375_gl_ram_n_552, FE_PHN374_ml_il_color1_n_10, FE_PHN373_ml_ms_cnt_n_21 : std_logic;
  signal FE_PHN372_ml_ms_n_57, FE_PHN371_gl_vgd_n_64, FE_PHN370_gl_ram_n_243, FE_PHN369_gl_ram_n_237, FE_PHN368_ml_ms_cnt_n_22 : std_logic;
  signal FE_PHN367_ml_ms_mfsm_n_36, FE_PHN366_gl_ram_n_568, FE_PHN365_gl_ram_n_80, FE_PHN364_gl_gr_lg_lv_n_14, FE_PHN363_ml_ms_cnt_n_19 : std_logic;
  signal FE_PHN362_gl_sig_v, FE_PHN361_gl_ram_n_78, FE_PHN360_gl_ram_n_142, FE_PHN359_gl_ram_n_77, FE_PHN358_gl_sig_scale_v : std_logic;
  signal FE_PHN357_gl_sig_scale_h, FE_PHN356_gl_gr_lg_sig_countdown_10, FE_PHN355_gl_gr_lg_sig_countdown_5, FE_PHN354_gl_gr_lg_sig_countdown_2, FE_PHN353_gl_gr_lg_sig_countdown_0 : std_logic;
  signal FE_PHN352_gl_gr_lg_sig_countdown_1, FE_PHN351_sig_logic_x_0, FE_PHN350_ml_ms_mfsm_state_4, FE_PHN349_sig_logic_y_0, FE_PHN348_gl_gr_lg_local_y_0 : std_logic;
  signal FE_PHN347_ml_ms_mfsm_state_3, FE_PHN346_gl_vgd_horizontal_counter_4, FE_PHN345_gl_vgd_horizontal_counter_1, FE_PHN344_gl_vgd_horizontal_counter_2, FE_PHN343_gl_vgd_horizontal_counter_5 : std_logic;
  signal FE_PHN342_gl_vgd_horizontal_counter_3, FE_PHN341_ml_ms_cnt_count_1, FE_PHN340_gl_vgd_horizontal_counter_0, FE_PHN339_gl_vgd_horizontal_counter_9, FE_PHN338_ml_ms_mfsm_state_2 : std_logic;
  signal FE_PHN337_gl_vgd_vertical_counter_2, FE_PHN336_gl_vgd_vertical_counter_0, FE_PHN335_ml_ms_count15k_1, FE_PHN334_ml_ms_count15k_0, FE_PHN333_gl_vgd_vertical_counter_1 : std_logic;
  signal FE_PHN332_ml_ms_count25M_8, FE_PHN331_gl_vgd_vertical_counter_9, FE_PHN330_gl_vgd_vertical_counter_6, FE_PHN329_ml_ms_mfsm_n_53, FE_PHN328_gl_vgd_vertical_counter_7 : std_logic;
  signal FE_PHN327_gl_ram_n_5, FE_PHN326_gl_vgd_vertical_counter_5, FE_PHN325_gl_gr_lg_lv_sig_edges, FE_PHN324_gl_vgd_vertical_counter_4, FE_PHN323_ml_ms_count25M_9 : std_logic;
  signal FE_PHN322_gl_vgd_vertical_counter_3, FE_PHN321_gl_vgd_n_77, FE_PHN320_ml_buttons_mouse_3, FE_PHN319_gl_gr_lg_sig_countdown_3, FE_PHN318_ml_ms_count25M_6 : std_logic;
  signal FE_PHN317_gl_ram_ram_86_1, FE_PHN316_gl_ram_ram_10_0, FE_PHN315_gl_ram_ram_61_1, FE_PHN314_gl_ram_ram_46_2, FE_PHN313_ml_ms_cntD_count_1 : std_logic;
  signal FE_PHN312_gl_ram_ram_80_0, FE_PHN311_gl_ram_ram_5_0, FE_PHN310_gl_ram_ram_20_2, FE_PHN309_gl_ram_ram_37_0, FE_PHN308_ml_ms_count25M_5 : std_logic;
  signal FE_PHN307_data_in, FE_PHN306_gl_ram_ram_39_2, FE_PHN305_gl_ram_ram_70_2, FE_PHN304_gl_gr_lg_lcountdown_l_edge_reg1, FE_PHN303_gl_ram_ram_71_1 : std_logic;
  signal FE_PHN302_gl_ram_ram_87_2, FE_PHN301_gl_gr_lg_lh_n_21, FE_PHN300_gl_gr_lg_lh_n_14, FE_PHN299_ml_ms_data_sr_11bit_7, FE_PHN298_gl_ram_ram_86_2 : std_logic;
  signal FE_PHN297_gl_Hint, FE_PHN296_gl_ram_ram_78_1, FE_PHN295_gl_ram_ram_14_2, FE_PHN294_gl_ram_ram_82_2, FE_PHN293_gl_ram_ram_39_0 : std_logic;
  signal FE_PHN292_gl_ram_ram_14_0, FE_PHN291_gl_ram_ram_86_0, FE_PHN290_gl_ram_ram_53_0, FE_PHN289_gl_ram_ram_46_1, FE_PHN288_gl_ram_ram_38_1 : std_logic;
  signal FE_PHN287_gl_ram_ram_23_2, FE_PHN286_gl_ram_ram_76_0, FE_PHN285_gl_ram_ram_36_1, FE_PHN284_ml_mouseY_0, FE_PHN283_gl_ram_ram_53_1 : std_logic;
  signal FE_PHN282_gl_ram_ram_23_1, FE_PHN281_gl_ram_ram_22_1, FE_PHN280_gl_ram_ram_66_2, FE_PHN279_ml_ms_data_sr_11bit_2, FE_PHN278_gl_ram_ram_52_2 : std_logic;
  signal FE_PHN277_gl_ram_ram_63_1, FE_PHN276_gl_ram_ram_55_1, FE_PHN275_ml_ms_data_sr_11bit_3, FE_PHN274_gl_ram_ram_36_0, FE_PHN273_gl_ram_ram_63_0 : std_logic;
  signal FE_PHN272_gl_ram_ram_47_0, FE_PHN271_gl_ram_ram_87_1, FE_PHN270_gl_ram_ram_76_2, FE_PHN269_gl_ram_ram_6_0, FE_PHN268_gl_ram_ram_6_1 : std_logic;
  signal FE_PHN267_gl_ram_ram_15_2, FE_PHN266_gl_ram_ram_13_0, FE_PHN265_gl_ram_ram_22_0, FE_PHN264_gl_ram_ram_68_0, FE_PHN263_gl_ram_ram_6_2 : std_logic;
  signal FE_PHN262_gl_ram_ram_55_2, FE_PHN261_gl_ram_ram_54_1, FE_PHN260_gl_ram_ram_45_1, FE_PHN259_gl_ram_ram_95_2, FE_PHN258_gl_ram_ram_30_1 : std_logic;
  signal FE_PHN257_gl_ram_ram_98_0, FE_PHN256_gl_ram_ram_99_0, FE_PHN255_gl_ram_ram_70_0, FE_PHN254_gl_ram_ram_63_2, FE_PHN253_gl_ram_ram_61_0 : std_logic;
  signal FE_PHN252_gl_ram_ram_64_2, FE_PHN251_gl_ram_ram_28_0, FE_PHN250_gl_ram_ram_69_2, FE_PHN249_gl_ram_ram_55_0, FE_PHN248_gl_ram_ram_99_1 : std_logic;
  signal FE_PHN247_gl_ram_ram_58_2, FE_PHN246_gl_ram_ram_74_1, FE_PHN245_gl_ram_ram_20_0, FE_PHN244_gl_ram_ram_61_2, FE_PHN243_gl_ram_ram_4_1 : std_logic;
  signal FE_PHN242_gl_ram_ram_81_2, FE_PHN241_gl_ram_ram_90_2, FE_PHN240_gl_ram_ram_78_2, FE_PHN239_gl_ram_ram_34_2, FE_PHN238_gl_ram_ram_79_2 : std_logic;
  signal FE_PHN237_gl_ram_ram_29_2, FE_PHN236_gl_ram_ram_85_1, FE_PHN235_gl_ram_ram_89_2, FE_PHN234_gl_ram_ram_74_2, FE_PHN233_gl_ram_ram_94_0 : std_logic;
  signal FE_PHN232_gl_ram_ram_62_1, FE_PHN231_gl_ram_ram_47_1, FE_PHN230_gl_ram_ram_84_1, FE_PHN229_gl_ram_ram_69_1, FE_PHN228_gl_ram_ram_59_0 : std_logic;
  signal FE_PHN227_gl_ram_ram_49_1, FE_PHN226_gl_ram_ram_77_2, FE_PHN225_gl_ram_ram_44_2, FE_PHN224_gl_ram_ram_95_1, FE_PHN223_gl_ram_ram_26_1 : std_logic;
  signal FE_PHN222_gl_ram_ram_41_1, FE_PHN221_gl_ram_ram_64_0, FE_PHN220_gl_ram_ram_93_0, FE_PHN219_gl_ram_ram_81_1, FE_PHN218_gl_ram_ram_26_2 : std_logic;
  signal FE_PHN217_gl_ram_ram_32_2, FE_PHN216_gl_ram_ram_89_1, FE_PHN215_gl_ram_ram_69_0, FE_PHN214_gl_ram_ram_98_1, FE_PHN213_gl_ram_ram_49_0 : std_logic;
  signal FE_PHN212_gl_ram_ram_75_1, FE_PHN211_gl_ram_ram_57_0, FE_PHN210_gl_ram_ram_96_0, FE_PHN209_gl_ram_ram_80_2, FE_PHN208_gl_ram_ram_49_2 : std_logic;
  signal FE_PHN207_gl_ram_ram_62_2, FE_PHN206_gl_ram_ram_47_2, FE_PHN205_gl_ram_ram_14_1, FE_PHN204_gl_ram_ram_15_0, FE_PHN203_gl_ram_ram_2_1 : std_logic;
  signal FE_PHN202_gl_ram_ram_38_2, FE_PHN201_gl_ram_ram_30_0, FE_PHN200_gl_ram_ram_67_1, FE_PHN199_gl_ram_ram_77_1, FE_PHN198_gl_ram_ram_54_2 : std_logic;
  signal FE_PHN197_ml_il_y1_state_0, FE_PHN196_gl_ram_ram_72_2, FE_PHN195_gl_ram_ram_7_0, FE_PHN194_gl_ram_ram_1_1, FE_PHN193_gl_ram_ram_90_1 : std_logic;
  signal FE_PHN192_gl_ram_ram_16_0, FE_PHN191_gl_ram_ram_75_2, FE_PHN190_gl_ram_ram_93_1, FE_PHN189_gl_ram_ram_76_1, FE_PHN188_gl_ram_ram_83_2 : std_logic;
  signal FE_PHN187_gl_ram_ram_34_0, FE_PHN186_gl_ram_ram_30_2, FE_PHN185_gl_ram_ram_58_0, FE_PHN184_gl_ram_ram_21_1, FE_PHN183_gl_ram_ram_22_2 : std_logic;
  signal FE_PHN182_gl_ram_ram_25_2, FE_PHN181_gl_gr_lg_lh_n_17, FE_PHN180_gl_ram_ram_39_1, FE_PHN179_gl_ram_ram_51_0, FE_PHN178_gl_ram_ram_52_0 : std_logic;
  signal FE_PHN177_gl_ram_ram_13_2, FE_PHN176_gl_ram_ram_26_0, FE_PHN175_gl_ram_ram_15_1, FE_PHN174_gl_ram_ram_31_1, FE_PHN173_gl_ram_ram_7_1 : std_logic;
  signal FE_PHN172_gl_ram_ram_31_0, FE_PHN171_gl_ram_ram_3_1, FE_PHN170_ml_il_x1_state_0, FE_PHN169_gl_ram_ram_35_1, FE_PHN168_gl_ram_ram_91_0 : std_logic;
  signal FE_PHN167_gl_ram_ram_42_0, FE_PHN166_gl_ram_ram_10_2, FE_PHN165_gl_ram_ram_48_0, FE_PHN164_gl_ram_ram_91_2, FE_PHN163_gl_ram_ram_40_2 : std_logic;
  signal FE_PHN162_gl_ram_ram_74_0, FE_PHN161_gl_ram_ram_85_0, FE_PHN160_gl_ram_ram_10_1, FE_PHN159_gl_ram_ram_92_0, FE_PHN158_gl_ram_ram_19_2 : std_logic;
  signal FE_PHN157_gl_ram_ram_70_1, FE_PHN156_gl_ram_ram_94_2, FE_PHN155_gl_ram_ram_23_0, FE_PHN154_gl_ram_ram_84_0, FE_PHN153_gl_ram_ram_83_1 : std_logic;
  signal FE_PHN152_gl_ram_ram_79_0, FE_PHN151_gl_ram_ram_28_2, FE_PHN150_gl_ram_ram_81_0, FE_PHN149_gl_ram_ram_9_1, FE_PHN148_gl_ram_ram_56_0 : std_logic;
  signal FE_PHN147_gl_ram_ram_90_0, FE_PHN146_gl_ram_ram_38_0, FE_PHN145_gl_ram_ram_45_2, FE_PHN144_gl_ram_ram_65_1, FE_PHN143_gl_ram_ram_66_1 : std_logic;
  signal FE_PHN142_gl_ram_ram_93_2, FE_PHN141_gl_ram_ram_78_0, FE_PHN140_gl_ram_ram_12_0, FE_PHN139_gl_ram_ram_72_1, FE_PHN138_gl_ram_ram_46_0 : std_logic;
  signal FE_PHN137_gl_ram_ram_28_1, FE_PHN136_gl_ram_ram_18_1, FE_PHN135_gl_ram_ram_79_1, FE_PHN134_gl_ram_ram_57_2, FE_PHN133_gl_ram_ram_52_1 : std_logic;
  signal FE_PHN132_gl_ram_ram_80_1, FE_PHN131_gl_ram_ram_17_0, FE_PHN130_gl_ram_ram_71_0, FE_PHN129_gl_ram_ram_71_2, FE_PHN128_gl_ram_ram_68_1 : std_logic;
  signal FE_PHN127_gl_ram_ram_37_1, FE_PHN126_gl_ram_ram_13_1, FE_PHN125_gl_ram_ram_65_0, FE_PHN124_gl_ram_ram_62_0, FE_PHN123_ml_ms_count_debounce_11 : std_logic;
  signal FE_PHN122_gl_ram_ram_51_1, FE_PHN121_gl_ram_ram_50_0, FE_PHN120_gl_ram_ram_45_0, FE_PHN119_gl_ram_ram_29_0, FE_PHN118_gl_ram_ram_59_1 : std_logic;
  signal FE_PHN117_gl_ram_ram_53_2, FE_PHN116_gl_ram_ram_67_2, FE_PHN115_gl_ram_ram_95_0, FE_PHN114_gl_ram_ram_64_1, FE_PHN113_gl_ram_ram_99_2 : std_logic;
  signal FE_PHN112_gl_ram_ram_87_0, FE_PHN111_gl_ram_ram_44_1, FE_PHN110_gl_ram_ram_88_2, FE_PHN109_gl_ram_ram_85_2, FE_PHN108_gl_ram_ram_92_2 : std_logic;
  signal FE_PHN107_gl_ram_ram_72_0, FE_PHN106_gl_ram_ram_94_1, FE_PHN105_gl_ram_ram_21_2, FE_PHN104_gl_ram_ram_88_1, FE_PHN103_gl_ram_ram_68_2 : std_logic;
  signal FE_PHN102_gl_ram_ram_5_2, FE_PHN101_gl_ram_ram_92_1, FE_PHN100_gl_ram_ram_54_0, FE_PHN99_gl_ram_ram_97_2, FE_PHN98_gl_ram_ram_77_0 : std_logic;
  signal FE_PHN97_gl_ram_ram_16_1, FE_PHN96_gl_ram_ram_17_2, FE_PHN95_gl_ram_ram_7_2, FE_PHN94_gl_ram_ram_4_2, FE_PHN93_gl_gr_lg_lh_n_15 : std_logic;
  signal FE_PHN92_gl_ram_ram_84_2, FE_PHN91_ml_ms_cnt_n_0, FE_PHN90_ml_ms_data_sr_11bit_4, FE_PHN89_ml_ms_cntD_n_0, FE_PHN88_gl_vga_buf_Vint : std_logic;
  signal FE_PHN87_ml_il_color1_state_hs_0, FE_PHN86_ml_ms_sr11_data_out_0_79, FE_PHN85_ml_mouseX_2, FE_PHN84_ml_mouseX_1, FE_PHN83_clk15k_in : std_logic;
  signal FE_PHN82_ml_mouseY_2, FE_PHN81_gl_vga_buf_Bint, FE_PHN80_ml_ms_sr11_data_out_5_84, FE_PHN79_ml_mouseY_1, FE_PHN78_ml_ms_sr11_data_out_1_80 : std_logic;
  signal FE_PHN77_ml_ms_n_26, FE_PHN76_ml_mouseX_0, FE_PHN75_ml_ms_n_20, FE_PHN74_ml_ms_n_19, FE_PHN73_ml_ms_n_25 : std_logic;
  signal FE_PHN72_ml_ms_data_sr_11bit_6, FE_PHN71_gl_vga_buf_Rint, FE_PHN70_gl_vga_buf_Hint, FE_PHN69_ml_ms_count_debounce_5, FE_PHN68_ml_ms_count_debounce_reset : std_logic;
  signal FE_PHN67_gl_vga_buf_Gint, FE_PHN66_gl_vgd_vertical_9, FE_PHN65_ml_ms_count_debounce_4, FE_PHN64_ml_ms_count_debounce_3, FE_PHN63_ml_ms_count25M_7 : std_logic;
  signal FE_PHN62_ml_ms_count_debounce_8, FE_PHN61_ml_ms_count_debounce_9, FE_PHN60_ml_ms_cntD_count_0, FE_PHN59_ml_il_color1_n_1, FE_PHN58_ml_ms_cntD_count_2 : std_logic;
  signal FE_PHN57_gl_vgd_vertical_counter_8, FE_PHN56_ml_il_x1_state_1, FE_PHN55_ml_buttons_mouse_4, FE_PHN54_ml_il_y1_state_1, FE_PHN53_ml_ms_ed_reg1 : std_logic;
  signal FE_PHN52_gl_gr_lg_lv_l_edge_reg1, FE_PHN51_gl_gr_lg_lh_l_edge_reg1, FE_PHN50_gl_gr_lg_le_new_count_e_0, FE_PHN49_gl_gr_lg_le_new_count_e_1, FE_PHN48_gl_gr_lg_le_new_count_e_7 : std_logic;
  signal FE_PHN47_gl_gr_lg_le_new_count_e_2, FE_PHN46_gl_gr_lg_le_new_count_e_4, FE_PHN45_gl_gr_lg_le_new_count_e_9, FE_PHN44_gl_gr_lg_le_new_count_e_3, FE_PHN43_gl_gr_lg_le_new_count_e_8 : std_logic;
  signal FE_PHN42_gl_gr_lg_le_new_count_e_5, FE_PHN41_gl_gr_lg_le_new_count_e_6, FE_OFN40_gl_ram_n_16, FE_OFN39_gl_ram_n_16, FE_OFN38_gl_ram_n_16 : std_logic;
  signal FE_OFN37_gl_ram_n_16, FE_OFN36_clk15k_switch, FE_OFN35_reset, FE_OFN34_R, FE_OFN33_B : std_logic;
  signal FE_OFN32_G, FE_OFN31_H, FE_OFN30_V, FE_OFN29_gl_rom_n_20, FE_OFN28_gl_rom_n_20 : std_logic;
  signal FE_OFN27_gl_rom_n_20, FE_OFN26_gl_rom_n_19, FE_OFN25_gl_rom_n_19, FE_OFN24_gl_rom_n_19, FE_OFN23_gl_rom_n_21 : std_logic;
  signal FE_OFN22_gl_rom_n_21, FE_OFN21_gl_rom_n_21, FE_OFN20_gl_rom_n_21, FE_OFN19_gl_rom_n_21, FE_OFN18_gl_rom_n_15 : std_logic;
  signal FE_OFN17_gl_rom_n_15, FE_OFN16_gl_rom_n_15, FE_OFN15_gl_rom_n_15, FE_OFN14_gl_rom_n_15, FE_OFN13_gl_rom_n_22 : std_logic;
  signal FE_OFN12_gl_rom_n_22, FE_OFN11_gl_rom_n_22, FE_OFN10_gl_rom_n_17, FE_OFN9_gl_rom_n_17, FE_OFN8_gl_rom_n_17 : std_logic;
  signal FE_OFN7_gl_rom_n_18, FE_OFN6_gl_rom_n_18, FE_OFN5_gl_rom_n_18, FE_OFN4_gl_rom_n_16, FE_OFN3_gl_rom_n_16 : std_logic;
  signal FE_OFN2_gl_rom_n_16, FE_OFN1_gl_rom_n_16, FE_OFN0_gl_rom_n_16, CTS_24, CTS_23 : std_logic;
  signal CTS_22, CTS_21, CTS_20, CTS_19, FE_DBTN0_reset : std_logic;
  signal ml_il_x1_input_register : std_logic_vector(3 downto 0);
  signal ml_mouseX : std_logic_vector(2 downto 0);
  signal sig_logic_x : std_logic_vector(3 downto 0);
  signal ml_buttons_mouse : std_logic_vector(4 downto 0);
  signal ml_il_x1_state : std_logic_vector(1 downto 0);
  signal ml_il_y1_input_register : std_logic_vector(3 downto 0);
  signal ml_mouseY : std_logic_vector(2 downto 0);
  signal sig_logic_y : std_logic_vector(3 downto 0);
  signal ml_il_y1_state : std_logic_vector(1 downto 0);
  signal gl_sig_x : std_logic_vector(3 downto 0);
  signal gl_sig_y : std_logic_vector(3 downto 0);
  signal gl_sig_rom : std_logic_vector(1 downto 0);
  signal gl_gr_lg_local_x : std_logic_vector(3 downto 0);
  signal gl_gr_lg_local_y : std_logic_vector(3 downto 0);
  signal sig_output_color : std_logic_vector(2 downto 0);
  signal gl_sig_ram : std_logic_vector(2 downto 0);
  signal gl_sig_e : std_logic_vector(9 downto 0);
  signal gl_rom_rom_776 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_779 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_385 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_389 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_977 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_981 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_980 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_982 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_384 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_387 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_978 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_979 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_976 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_983 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_712 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_713 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_956 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_958 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_882 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_887 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_706 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_711 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_985 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_989 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_988 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_990 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_378 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_383 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_986 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_987 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_984 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_991 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_708 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_710 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_380 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_382 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_994 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_999 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_993 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_997 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_880 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_883 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_381 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_379 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_996 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_998 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_376 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_377 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_992 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_995 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1020 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1023 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_709 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_707 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1018 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1022 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_362 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_367 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_704 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_705 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1017 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1021 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1016 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1019 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_361 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_365 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1004 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1007 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1002 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1006 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_364 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_366 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_360 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_363 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1001 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1005 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1000 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1003 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_972 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_975 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_957 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_955 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_970 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_974 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_370 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_375 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_969 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_973 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_852 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_855 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_968 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_971 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_372 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_374 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_794 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_799 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_964 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_967 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_373 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_371 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_962 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_966 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_850 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_854 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_961 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_965 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_960 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_963 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_368 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_369 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_953 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_793 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_797 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_796 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_798 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_338 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_343 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_954 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_340 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_342 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_952 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_959 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_792 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_795 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_937 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_941 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_341 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_339 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_940 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_942 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_938 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_939 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_336 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_337 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_936 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_943 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_924 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_927 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_849 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_853 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_922 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_926 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_346 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_351 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_921 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_925 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_806 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_805 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_920 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_923 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_348 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_350 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_848 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_851 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_930 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_935 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_929 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_933 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_349 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_347 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_932 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_934 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_344 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_345 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_928 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_931 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_804 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_801 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_945 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_949 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_948 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_950 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_354 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_359 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_802 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_807 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_946 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_947 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_356 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_358 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_944 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_951 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_914 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_919 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_800 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_803 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_357 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_355 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_913 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_917 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_352 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_353 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_918 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_915 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_912 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_916 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_910 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_909 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_908 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_905 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_329 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_333 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_906 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_911 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_904 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_907 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_332 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_334 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_817 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_821 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_898 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_903 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_890 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_895 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_330 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_331 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_897 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_901 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_820 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_822 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_328 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_335 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_900 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_902 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_896 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_899 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_892 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_894 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_700 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_703 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_322 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_327 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_698 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_702 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_818 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_819 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_697 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_701 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_696 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_699 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_324 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_326 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_325 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_323 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_684 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_687 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_816 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_823 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_682 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_686 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_320 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_321 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_681 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_685 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_680 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_683 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_893 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_891 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_690 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_695 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_692 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_694 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_124 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_127 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_693 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_691 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_688 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_689 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_122 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_126 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_660 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_663 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_786 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_791 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_658 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_662 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_785 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_789 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_121 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_125 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_120 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_123 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_657 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_661 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_656 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_659 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_666 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_671 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_888 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_889 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_790 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_787 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_665 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_669 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_106 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_111 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_105 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_109 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_670 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_667 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_664 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_668 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_676 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_679 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_784 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_788 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_110 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_107 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_674 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_678 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_104 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_108 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_673 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_677 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_672 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_675 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_652 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_655 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_650 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_654 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_874 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_879 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_114 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_119 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_649 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_653 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_116 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_118 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_648 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_651 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_825 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_829 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_828 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_830 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_642 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_647 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_117 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_115 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_641 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_645 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_644 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_646 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_640 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_643 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_569 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_573 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_112 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_113 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_873 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_877 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_82 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_87 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_572 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_574 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_826 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_827 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_570 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_571 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_84 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_86 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_568 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_575 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_824 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_831 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_85 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_83 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_554 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_559 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_553 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_557 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_556 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_558 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_80 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_81 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_552 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_555 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_878 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_875 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_564 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_567 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_562 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_566 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_90 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_95 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_810 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_815 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_561 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_565 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_92 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_94 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_560 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_563 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_532 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_535 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_93 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_91 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_530 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_534 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_809 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_813 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_529 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_533 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_528 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_531 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_88 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_89 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_540 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_543 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_872 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_876 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_814 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_811 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_100 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_103 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_538 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_542 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_98 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_102 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_537 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_541 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_536 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_539 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_548 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_551 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_808 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_812 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_97 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_101 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_546 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_550 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_96 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_99 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_545 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_549 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_544 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_547 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_524 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_527 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_522 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_526 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_74 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_79 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_842 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_847 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_521 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_525 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_778 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_783 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_520 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_523 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_73 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_77 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_518 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_517 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_78 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_75 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_516 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_513 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_72 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_76 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_514 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_519 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_512 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_515 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_777 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_781 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_66 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_71 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_780 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_782 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_498 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_503 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_497 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_501 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_841 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_845 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_68 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_70 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_500 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_502 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_496 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_499 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_69 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_67 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1008 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1011 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_470 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_469 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_468 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_465 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_64 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_65 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_466 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_471 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_464 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_467 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_846 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_843 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_474 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_479 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_770 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_775 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_476 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_478 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_217 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_221 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_477 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_475 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_472 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_473 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_220 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_222 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_769 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_773 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_484 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_487 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_482 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_486 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_218 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_219 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_481 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_485 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_480 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_483 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_216 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_223 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_506 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_511 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_840 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_844 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_772 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_774 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_225 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_229 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_508 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_510 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_768 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_771 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_509 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_507 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_228 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_230 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_504 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_505 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_494 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_493 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_226 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_227 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_492 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_489 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1012 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1014 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_490 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_495 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_224 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_231 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_488 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_491 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_834 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_839 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_458 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_463 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_457 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_461 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_242 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_247 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_460 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_462 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_456 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_459 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_241 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_245 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_454 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_453 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_244 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_246 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_452 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_449 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_450 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_455 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_240 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_243 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_448 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_451 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_833 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_837 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_442 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_447 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_212 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_215 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_444 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_446 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_210 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_214 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_445 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_443 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_440 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_441 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_426 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_431 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_209 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_213 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_425 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_429 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_428 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_430 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_424 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_427 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_208 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_211 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_838 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_835 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_410 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_415 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_409 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_413 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_252 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_255 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_412 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_414 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_250 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_254 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_408 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_411 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_832 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_836 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_420 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_423 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_249 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_253 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_418 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_422 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_417 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_421 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_416 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_419 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_248 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_251 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_438 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_437 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_436 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_433 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_233 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_237 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_434 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_439 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_236 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_238 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_432 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_435 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_402 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_407 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_234 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_235 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_401 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_405 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_404 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_406 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_232 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_239 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_400 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_403 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_398 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_397 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_396 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_393 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_201 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_205 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_394 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_399 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_204 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_206 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_392 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_395 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_388 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_391 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_634 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_639 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_386 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_390 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_202 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_203 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_200 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_207 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_193 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_197 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_196 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_198 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_636 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_638 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_194 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_195 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_192 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_199 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_637 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_635 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_316 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_319 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_314 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_318 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_313 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_317 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_312 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_315 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_300 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_303 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_632 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_633 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_298 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_302 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_297 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_301 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_296 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_299 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_281 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_285 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_284 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_286 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_282 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_283 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_617 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_621 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_280 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_287 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_620 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_622 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_289 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_293 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_292 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_294 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_290 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_291 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_288 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_295 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_618 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_619 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_308 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_311 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_306 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_310 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_305 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_309 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_304 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_307 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_274 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_279 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_273 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_277 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_276 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_278 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_272 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_275 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_616 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_623 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_268 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_271 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_266 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_270 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_265 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_269 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_264 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_267 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_602 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_607 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_258 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_263 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_257 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_261 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_260 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_262 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_256 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_259 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_604 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_606 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_605 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_603 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_188 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_191 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_186 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_190 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_185 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_189 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_184 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_187 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_600 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_601 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_169 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_173 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_172 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_174 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_170 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_171 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_168 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_175 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_154 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_159 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_610 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_615 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_156 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_158 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_157 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_155 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_152 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_153 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_609 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_613 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_164 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_167 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_162 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_166 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_161 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_165 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_160 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_163 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_614 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_611 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_178 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_183 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_608 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_612 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_180 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_182 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_181 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_179 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_176 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_177 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_146 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_151 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_148 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_150 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_149 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_147 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_144 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_145 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_138 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_143 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_625 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_629 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_140 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_142 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_141 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_139 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_136 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_137 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_130 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_135 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_628 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_630 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_129 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_133 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_132 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_134 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_128 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_131 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_626 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_627 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_58 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_63 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_57 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_61 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_60 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_62 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_56 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_59 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_624 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_631 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_44 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_47 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_42 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_46 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_41 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_45 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_40 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_43 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1013 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_594 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_599 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_50 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_55 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_52 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_54 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_53 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_51 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_48 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_49 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_593 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_597 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_17 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_21 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_20 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_22 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_18 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_19 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_16 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_23 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_596 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_598 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_26 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_31 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_25 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_29 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_30 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_27 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_592 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_595 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_24 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_28 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_34 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_39 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_36 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_38 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_37 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_35 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_33 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_32 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_9 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_13 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_12 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_15 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_14 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_10 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_11 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_586 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_591 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_8 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_2 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_7 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_5 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_588 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_590 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_4 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_6 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_0 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_3 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_589 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_587 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_584 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_585 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_578 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_583 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_580 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_582 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_860 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_863 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_858 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_862 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_857 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_861 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_856 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_859 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_868 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_871 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_866 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_870 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_581 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_579 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_865 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_869 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_864 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_867 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_884 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_886 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_576 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_577 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_881 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_885 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_754 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_759 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_753 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_757 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_758 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_755 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_752 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_756 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_722 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_727 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_724 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_726 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1009 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_725 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_723 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_720 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_721 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_730 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_735 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_729 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_733 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_766 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_765 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_734 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_731 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_764 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_761 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_762 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_767 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_760 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_763 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_728 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_732 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_746 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_751 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_748 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_750 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_749 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_747 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_744 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_745 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_738 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_743 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_740 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_742 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_741 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_739 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_736 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_737 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_714 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_719 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_716 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_718 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_717 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_715 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1010 : std_logic_vector(1 downto 0);
  signal gl_rom_rom_1015 : std_logic_vector(1 downto 0);
  signal gl_ram_ram_96 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_97 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_98 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_99 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_88 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_91 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_41 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_42 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_62 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_63 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_60 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_61 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_44 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_45 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_57 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_58 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_40 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_43 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_56 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_59 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_72 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_75 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_54 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_55 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_49 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_50 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_52 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_53 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_38 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_39 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_48 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_51 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_33 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_34 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_30 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_31 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_24 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_27 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_36 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_37 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_28 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_29 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_86 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_87 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_25 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_26 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_32 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_35 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_14 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_15 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_12 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_13 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_66 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_67 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_10 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_11 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_80 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_83 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_8 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_9 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_46 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_47 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_84 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_85 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_78 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_79 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_81 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_82 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_22 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_23 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_16 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_19 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_20 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_21 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_17 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_18 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_70 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_71 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_6 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_7 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_1 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_2 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_4 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_5 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_0 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_3 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_94 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_95 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_65 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_68 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_69 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_92 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_93 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_89 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_90 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_64 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_73 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_74 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_76 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_77 : std_logic_vector(2 downto 0);
  signal gl_ram_ram_position : std_logic_vector(6 downto 0);
  signal gl_ram_x_grid : std_logic_vector(6 downto 0);
  signal gl_ram_y_grid : std_logic_vector(6 downto 0);
  signal gl_gr_lg_sig_countdown : std_logic_vector(10 downto 0);
  signal gl_gr_lg_le_new_count_e : std_logic_vector(9 downto 0);
  signal ml_ms_sfsm_state : std_logic_vector(3 downto 0);
  signal ml_ms_sr_new_new_data : std_logic_vector(8 downto 0);
  signal ml_ms_count25M : std_logic_vector(12 downto 0);
  signal ml_ms_data_sr_11bit : std_logic_vector(10 downto 0);
  signal ml_ms_btns : std_logic_vector(4 downto 0);
  signal ml_ms_mouse_x : std_logic_vector(2 downto 0);
  signal ml_ms_mouse_y : std_logic_vector(2 downto 0);
  signal ml_ms_mfsm_state : std_logic_vector(4 downto 0);
  signal ml_ms_count15k : std_logic_vector(3 downto 0);
  signal ml_ms_cnt_count : std_logic_vector(12 downto 0);
  signal ml_ms_count_debounce : std_logic_vector(12 downto 0);
  signal ml_ms_cntD_count : std_logic_vector(12 downto 0);
  signal ml_il_color1_state : std_logic_vector(2 downto 0);
  signal ml_il_color1_state_hs : std_logic_vector(1 downto 0);
  signal gl_vgd_horizontal : std_logic_vector(9 downto 0);
  signal gl_vgd_vertical : std_logic_vector(9 downto 0);
  signal gl_vgd_horizontal_counter : std_logic_vector(9 downto 0);
  signal gl_vgd_vertical_counter : std_logic_vector(9 downto 0);
  signal ml_ms_ed_state : std_logic_vector(1 downto 0);
  signal UNCONNECTED, UNCONNECTED0, UNCONNECTED1, gl_Bint, gl_Gint : std_logic;
  signal gl_Hint, gl_Rint, gl_const_gr_lg_mul_88_58_n_1, gl_const_gr_lg_mul_88_58_n_3, gl_const_gr_lg_mul_88_58_n_4 : std_logic;
  signal gl_const_gr_lg_mul_88_58_n_5, gl_const_gr_lg_mul_88_58_n_6, gl_const_gr_lg_mul_88_58_n_7, gl_const_gr_lg_mul_88_58_n_8, gl_const_gr_lg_mul_88_58_n_9 : std_logic;
  signal gl_const_gr_lg_mul_88_58_n_10, gl_const_gr_lg_mul_88_58_n_11, gl_const_gr_lg_mul_88_58_n_12, gl_const_gr_lg_mul_88_58_n_13, gl_const_gr_lg_mul_88_58_n_14 : std_logic;
  signal gl_const_gr_lg_mul_88_58_n_15, gl_const_gr_lg_mul_88_58_n_16, gl_const_gr_lg_mul_88_58_n_17, gl_const_gr_lg_mul_88_58_n_18, gl_const_gr_lg_mul_88_58_n_19 : std_logic;
  signal gl_const_gr_lg_mul_88_58_n_20, gl_const_gr_lg_mul_88_58_n_21, gl_const_gr_lg_mul_88_58_n_22, gl_const_gr_lg_mul_88_58_n_23, gl_const_gr_lg_mul_88_58_n_25 : std_logic;
  signal gl_const_gr_lg_mul_88_58_n_27, gl_const_gr_lg_mul_88_58_n_29, gl_const_gr_lg_mul_88_58_n_31, gl_const_gr_lg_mul_88_58_n_33, gl_const_gr_lg_mul_88_58_n_35 : std_logic;
  signal gl_const_gr_lg_mul_88_58_n_37, gl_const_gr_lg_mul_88_58_n_39, gl_const_gr_lg_mul_88_58_n_41, gl_gr_lg_div_88_62_n_1, gl_gr_lg_div_88_62_n_2 : std_logic;
  signal gl_gr_lg_div_88_62_n_3, gl_gr_lg_div_88_62_n_4, gl_gr_lg_div_88_62_n_5, gl_gr_lg_div_88_62_n_6, gl_gr_lg_div_88_62_n_7 : std_logic;
  signal gl_gr_lg_div_88_62_n_8, gl_gr_lg_div_88_62_n_9, gl_gr_lg_div_88_62_n_10, gl_gr_lg_div_88_62_n_11, gl_gr_lg_div_88_62_n_12 : std_logic;
  signal gl_gr_lg_div_88_62_n_13, gl_gr_lg_div_88_62_n_14, gl_gr_lg_div_88_62_n_15, gl_gr_lg_div_88_62_n_16, gl_gr_lg_div_88_62_n_17 : std_logic;
  signal gl_gr_lg_div_88_62_n_18, gl_gr_lg_div_88_62_n_19, gl_gr_lg_div_88_62_n_20, gl_gr_lg_div_88_62_n_21, gl_gr_lg_div_88_62_n_22 : std_logic;
  signal gl_gr_lg_div_88_62_n_23, gl_gr_lg_div_88_62_n_24, gl_gr_lg_div_88_62_n_25, gl_gr_lg_div_88_62_n_26, gl_gr_lg_div_88_62_n_27 : std_logic;
  signal gl_gr_lg_div_88_62_n_28, gl_gr_lg_div_88_62_n_29, gl_gr_lg_div_88_62_n_30, gl_gr_lg_div_88_62_n_31, gl_gr_lg_div_88_62_n_32 : std_logic;
  signal gl_gr_lg_div_88_62_n_33, gl_gr_lg_div_88_62_n_34, gl_gr_lg_div_88_62_n_35, gl_gr_lg_div_88_62_n_36, gl_gr_lg_div_88_62_n_37 : std_logic;
  signal gl_gr_lg_div_88_62_n_38, gl_gr_lg_div_88_62_n_39, gl_gr_lg_div_88_62_n_40, gl_gr_lg_div_88_62_n_41, gl_gr_lg_div_88_62_n_42 : std_logic;
  signal gl_gr_lg_div_88_62_n_43, gl_gr_lg_div_88_62_n_44, gl_gr_lg_div_88_62_n_45, gl_gr_lg_div_88_62_n_46, gl_gr_lg_div_88_62_n_47 : std_logic;
  signal gl_gr_lg_div_88_62_n_48, gl_gr_lg_div_88_62_n_49, gl_gr_lg_div_88_62_n_50, gl_gr_lg_div_88_62_n_51, gl_gr_lg_div_88_62_n_52 : std_logic;
  signal gl_gr_lg_div_88_62_n_53, gl_gr_lg_div_88_62_n_54, gl_gr_lg_div_88_62_n_55, gl_gr_lg_div_88_62_n_56, gl_gr_lg_div_88_62_n_57 : std_logic;
  signal gl_gr_lg_div_88_62_n_58, gl_gr_lg_div_88_62_n_59, gl_gr_lg_div_88_62_n_60, gl_gr_lg_div_88_62_n_61, gl_gr_lg_div_88_62_n_62 : std_logic;
  signal gl_gr_lg_div_88_62_n_63, gl_gr_lg_div_88_62_n_64, gl_gr_lg_div_88_62_n_65, gl_gr_lg_div_88_62_n_66, gl_gr_lg_div_88_62_n_67 : std_logic;
  signal gl_gr_lg_div_88_62_n_68, gl_gr_lg_div_88_62_n_69, gl_gr_lg_div_88_62_n_70, gl_gr_lg_div_88_62_n_71, gl_gr_lg_div_88_62_n_73 : std_logic;
  signal gl_gr_lg_div_88_62_n_74, gl_gr_lg_div_88_62_n_75, gl_gr_lg_div_88_62_n_76, gl_gr_lg_div_88_62_n_77, gl_gr_lg_div_88_62_n_78 : std_logic;
  signal gl_gr_lg_div_88_62_n_79, gl_gr_lg_div_88_62_n_80, gl_gr_lg_div_88_62_n_81, gl_gr_lg_div_88_62_n_82, gl_gr_lg_div_88_62_n_83 : std_logic;
  signal gl_gr_lg_div_88_62_n_84, gl_gr_lg_div_88_62_n_85, gl_gr_lg_div_88_62_n_86, gl_gr_lg_div_88_62_n_87, gl_gr_lg_div_88_62_n_88 : std_logic;
  signal gl_gr_lg_div_88_62_n_89, gl_gr_lg_div_88_62_n_90, gl_gr_lg_div_88_62_n_91, gl_gr_lg_div_88_62_n_92, gl_gr_lg_div_88_62_n_93 : std_logic;
  signal gl_gr_lg_div_88_62_n_95, gl_gr_lg_div_88_62_n_96, gl_gr_lg_div_88_62_n_97, gl_gr_lg_div_88_62_n_99, gl_gr_lg_div_88_62_n_100 : std_logic;
  signal gl_gr_lg_div_88_62_n_101, gl_gr_lg_div_88_62_n_102, gl_gr_lg_div_88_62_n_103, gl_gr_lg_div_88_62_n_104, gl_gr_lg_div_88_62_n_105 : std_logic;
  signal gl_gr_lg_div_88_62_n_106, gl_gr_lg_div_88_62_n_107, gl_gr_lg_div_88_62_n_108, gl_gr_lg_div_88_62_n_109, gl_gr_lg_div_88_62_n_110 : std_logic;
  signal gl_gr_lg_div_88_62_n_111, gl_gr_lg_div_88_62_n_112, gl_gr_lg_div_88_62_n_113, gl_gr_lg_div_88_62_n_114, gl_gr_lg_div_88_62_n_115 : std_logic;
  signal gl_gr_lg_div_88_62_n_116, gl_gr_lg_div_88_62_n_117, gl_gr_lg_div_88_62_n_118, gl_gr_lg_div_88_62_n_119, gl_gr_lg_div_88_62_n_121 : std_logic;
  signal gl_gr_lg_div_88_62_n_122, gl_gr_lg_div_88_62_n_123, gl_gr_lg_div_88_62_n_125, gl_gr_lg_div_88_62_n_126, gl_gr_lg_div_88_62_n_127 : std_logic;
  signal gl_gr_lg_div_88_62_n_128, gl_gr_lg_div_88_62_n_129, gl_gr_lg_div_88_62_n_130, gl_gr_lg_div_88_62_n_131, gl_gr_lg_div_88_62_n_132 : std_logic;
  signal gl_gr_lg_div_88_62_n_133, gl_gr_lg_div_88_62_n_134, gl_gr_lg_div_88_62_n_135, gl_gr_lg_div_88_62_n_136, gl_gr_lg_div_88_62_n_137 : std_logic;
  signal gl_gr_lg_lcountdown_l_edge_reg1, gl_gr_lg_lcountdown_l_edge_reg2, gl_gr_lg_lcountdown_n_0, gl_gr_lg_lcountdown_n_1, gl_gr_lg_lcountdown_n_2 : std_logic;
  signal gl_gr_lg_lcountdown_n_3, gl_gr_lg_lcountdown_n_4, gl_gr_lg_lcountdown_n_5, gl_gr_lg_lcountdown_n_6, gl_gr_lg_lcountdown_n_7 : std_logic;
  signal gl_gr_lg_lcountdown_n_8, gl_gr_lg_lcountdown_n_9, gl_gr_lg_lcountdown_n_10, gl_gr_lg_lcountdown_n_11, gl_gr_lg_lcountdown_n_12 : std_logic;
  signal gl_gr_lg_lcountdown_n_13, gl_gr_lg_lcountdown_n_14, gl_gr_lg_lcountdown_n_15, gl_gr_lg_lcountdown_n_16, gl_gr_lg_lcountdown_n_17 : std_logic;
  signal gl_gr_lg_lcountdown_n_18, gl_gr_lg_lcountdown_n_19, gl_gr_lg_lcountdown_n_20, gl_gr_lg_lcountdown_n_21, gl_gr_lg_lcountdown_n_22 : std_logic;
  signal gl_gr_lg_lcountdown_n_23, gl_gr_lg_lcountdown_n_29, gl_gr_lg_lcountdown_sig_edge_fall, gl_gr_lg_le_n_0, gl_gr_lg_le_n_1 : std_logic;
  signal gl_gr_lg_le_n_2, gl_gr_lg_le_n_3, gl_gr_lg_le_n_4, gl_gr_lg_le_n_5, gl_gr_lg_le_n_6 : std_logic;
  signal gl_gr_lg_le_n_7, gl_gr_lg_le_n_8, gl_gr_lg_le_n_9, gl_gr_lg_le_n_10, gl_gr_lg_le_n_11 : std_logic;
  signal gl_gr_lg_le_n_12, gl_gr_lg_le_n_13, gl_gr_lg_le_n_14, gl_gr_lg_le_n_15, gl_gr_lg_le_n_16 : std_logic;
  signal gl_gr_lg_le_n_17, gl_gr_lg_le_n_18, gl_gr_lg_le_n_19, gl_gr_lg_le_n_20, gl_gr_lg_le_n_21 : std_logic;
  signal gl_gr_lg_le_n_22, gl_gr_lg_le_n_23, gl_gr_lg_le_n_24, gl_gr_lg_le_n_25, gl_gr_lg_le_n_26 : std_logic;
  signal gl_gr_lg_le_n_27, gl_gr_lg_le_n_28, gl_gr_lg_le_n_29, gl_gr_lg_le_n_31, gl_gr_lg_le_n_32 : std_logic;
  signal gl_gr_lg_lh_l_edge_n_0, gl_gr_lg_lh_l_edge_reg1, gl_gr_lg_lh_l_edge_reg2, gl_gr_lg_lh_n_3, gl_gr_lg_lh_n_4 : std_logic;
  signal gl_gr_lg_lh_n_5, gl_gr_lg_lh_n_6, gl_gr_lg_lh_n_7, gl_gr_lg_lh_n_8, gl_gr_lg_lh_n_10 : std_logic;
  signal gl_gr_lg_lh_n_12, gl_gr_lg_lh_n_13, gl_gr_lg_lh_n_14, gl_gr_lg_lh_n_15, gl_gr_lg_lh_n_16 : std_logic;
  signal gl_gr_lg_lh_n_17, gl_gr_lg_lh_n_21, gl_gr_lg_lh_sig_edges, gl_gr_lg_lv_l_edge_n_0, gl_gr_lg_lv_l_edge_reg1 : std_logic;
  signal gl_gr_lg_lv_l_edge_reg2, gl_gr_lg_lv_n_0, gl_gr_lg_lv_n_1, gl_gr_lg_lv_n_3, gl_gr_lg_lv_n_4 : std_logic;
  signal gl_gr_lg_lv_n_5, gl_gr_lg_lv_n_6, gl_gr_lg_lv_n_7, gl_gr_lg_lv_n_8, gl_gr_lg_lv_n_9 : std_logic;
  signal gl_gr_lg_lv_n_10, gl_gr_lg_lv_n_11, gl_gr_lg_lv_n_12, gl_gr_lg_lv_n_13, gl_gr_lg_lv_n_14 : std_logic;
  signal gl_gr_lg_lv_n_15, gl_gr_lg_lv_sig_edges, gl_gr_lg_n_104, gl_gr_lg_n_105, gl_gr_lg_n_113 : std_logic;
  signal gl_n_0, gl_n_1, gl_n_2, gl_n_3, gl_n_4 : std_logic;
  signal gl_n_5, gl_n_7, gl_n_8, gl_n_9, gl_n_10 : std_logic;
  signal gl_n_11, gl_n_12, gl_n_13, gl_n_14, gl_n_15 : std_logic;
  signal gl_n_16, gl_n_17, gl_n_19, gl_n_20, gl_n_21 : std_logic;
  signal gl_n_22, gl_n_23, gl_n_24, gl_n_25, gl_n_26 : std_logic;
  signal gl_n_27, gl_n_28, gl_n_29, gl_n_30, gl_n_31 : std_logic;
  signal gl_n_32, gl_n_33, gl_n_34, gl_n_35, gl_n_36 : std_logic;
  signal gl_n_37, gl_n_38, gl_n_39, gl_n_40, gl_n_41 : std_logic;
  signal gl_n_42, gl_n_43, gl_n_44, gl_n_45, gl_n_46 : std_logic;
  signal gl_n_47, gl_n_48, gl_n_49, gl_n_50, gl_n_51 : std_logic;
  signal gl_n_52, gl_n_53, gl_n_54, gl_n_55, gl_n_56 : std_logic;
  signal gl_n_57, gl_n_58, gl_n_59, gl_n_60, gl_n_61 : std_logic;
  signal gl_n_62, gl_n_63, gl_n_64, gl_n_65, gl_n_66 : std_logic;
  signal gl_n_84, gl_n_85, gl_n_86, gl_n_87, gl_n_88 : std_logic;
  signal gl_n_89, gl_n_90, gl_n_91, gl_n_92, gl_n_93 : std_logic;
  signal gl_n_94, gl_n_95, gl_n_96, gl_n_97, gl_n_98 : std_logic;
  signal gl_n_99, gl_n_100, gl_n_101, gl_n_102, gl_n_103 : std_logic;
  signal gl_n_125, gl_n_126, gl_ram_n_0, gl_ram_n_1, gl_ram_n_2 : std_logic;
  signal gl_ram_n_3, gl_ram_n_4, gl_ram_n_5, gl_ram_n_6, gl_ram_n_7 : std_logic;
  signal gl_ram_n_8, gl_ram_n_9, gl_ram_n_10, gl_ram_n_11, gl_ram_n_12 : std_logic;
  signal gl_ram_n_13, gl_ram_n_14, gl_ram_n_15, gl_ram_n_16, gl_ram_n_17 : std_logic;
  signal gl_ram_n_18, gl_ram_n_19, gl_ram_n_20, gl_ram_n_21, gl_ram_n_22 : std_logic;
  signal gl_ram_n_23, gl_ram_n_24, gl_ram_n_25, gl_ram_n_26, gl_ram_n_27 : std_logic;
  signal gl_ram_n_28, gl_ram_n_29, gl_ram_n_30, gl_ram_n_31, gl_ram_n_32 : std_logic;
  signal gl_ram_n_33, gl_ram_n_34, gl_ram_n_35, gl_ram_n_36, gl_ram_n_37 : std_logic;
  signal gl_ram_n_38, gl_ram_n_39, gl_ram_n_40, gl_ram_n_41, gl_ram_n_42 : std_logic;
  signal gl_ram_n_43, gl_ram_n_44, gl_ram_n_45, gl_ram_n_46, gl_ram_n_47 : std_logic;
  signal gl_ram_n_48, gl_ram_n_49, gl_ram_n_50, gl_ram_n_51, gl_ram_n_52 : std_logic;
  signal gl_ram_n_53, gl_ram_n_54, gl_ram_n_55, gl_ram_n_56, gl_ram_n_57 : std_logic;
  signal gl_ram_n_58, gl_ram_n_59, gl_ram_n_60, gl_ram_n_61, gl_ram_n_62 : std_logic;
  signal gl_ram_n_63, gl_ram_n_64, gl_ram_n_65, gl_ram_n_66, gl_ram_n_67 : std_logic;
  signal gl_ram_n_68, gl_ram_n_69, gl_ram_n_70, gl_ram_n_71, gl_ram_n_72 : std_logic;
  signal gl_ram_n_73, gl_ram_n_74, gl_ram_n_75, gl_ram_n_76, gl_ram_n_77 : std_logic;
  signal gl_ram_n_78, gl_ram_n_79, gl_ram_n_80, gl_ram_n_81, gl_ram_n_82 : std_logic;
  signal gl_ram_n_83, gl_ram_n_84, gl_ram_n_85, gl_ram_n_86, gl_ram_n_87 : std_logic;
  signal gl_ram_n_88, gl_ram_n_89, gl_ram_n_90, gl_ram_n_91, gl_ram_n_92 : std_logic;
  signal gl_ram_n_93, gl_ram_n_94, gl_ram_n_95, gl_ram_n_96, gl_ram_n_97 : std_logic;
  signal gl_ram_n_98, gl_ram_n_99, gl_ram_n_100, gl_ram_n_101, gl_ram_n_102 : std_logic;
  signal gl_ram_n_103, gl_ram_n_104, gl_ram_n_105, gl_ram_n_106, gl_ram_n_107 : std_logic;
  signal gl_ram_n_108, gl_ram_n_109, gl_ram_n_110, gl_ram_n_111, gl_ram_n_112 : std_logic;
  signal gl_ram_n_113, gl_ram_n_114, gl_ram_n_115, gl_ram_n_116, gl_ram_n_117 : std_logic;
  signal gl_ram_n_118, gl_ram_n_119, gl_ram_n_120, gl_ram_n_121, gl_ram_n_122 : std_logic;
  signal gl_ram_n_123, gl_ram_n_124, gl_ram_n_125, gl_ram_n_126, gl_ram_n_127 : std_logic;
  signal gl_ram_n_128, gl_ram_n_129, gl_ram_n_130, gl_ram_n_131, gl_ram_n_132 : std_logic;
  signal gl_ram_n_133, gl_ram_n_134, gl_ram_n_135, gl_ram_n_136, gl_ram_n_137 : std_logic;
  signal gl_ram_n_138, gl_ram_n_139, gl_ram_n_140, gl_ram_n_141, gl_ram_n_142 : std_logic;
  signal gl_ram_n_143, gl_ram_n_144, gl_ram_n_145, gl_ram_n_146, gl_ram_n_147 : std_logic;
  signal gl_ram_n_148, gl_ram_n_149, gl_ram_n_150, gl_ram_n_151, gl_ram_n_152 : std_logic;
  signal gl_ram_n_153, gl_ram_n_154, gl_ram_n_155, gl_ram_n_156, gl_ram_n_157 : std_logic;
  signal gl_ram_n_158, gl_ram_n_159, gl_ram_n_160, gl_ram_n_161, gl_ram_n_162 : std_logic;
  signal gl_ram_n_163, gl_ram_n_164, gl_ram_n_165, gl_ram_n_166, gl_ram_n_167 : std_logic;
  signal gl_ram_n_168, gl_ram_n_169, gl_ram_n_170, gl_ram_n_171, gl_ram_n_172 : std_logic;
  signal gl_ram_n_173, gl_ram_n_174, gl_ram_n_175, gl_ram_n_176, gl_ram_n_177 : std_logic;
  signal gl_ram_n_178, gl_ram_n_179, gl_ram_n_180, gl_ram_n_181, gl_ram_n_182 : std_logic;
  signal gl_ram_n_183, gl_ram_n_184, gl_ram_n_185, gl_ram_n_186, gl_ram_n_187 : std_logic;
  signal gl_ram_n_188, gl_ram_n_189, gl_ram_n_190, gl_ram_n_191, gl_ram_n_192 : std_logic;
  signal gl_ram_n_193, gl_ram_n_194, gl_ram_n_195, gl_ram_n_196, gl_ram_n_197 : std_logic;
  signal gl_ram_n_198, gl_ram_n_199, gl_ram_n_200, gl_ram_n_201, gl_ram_n_202 : std_logic;
  signal gl_ram_n_203, gl_ram_n_204, gl_ram_n_205, gl_ram_n_206, gl_ram_n_207 : std_logic;
  signal gl_ram_n_208, gl_ram_n_209, gl_ram_n_210, gl_ram_n_211, gl_ram_n_212 : std_logic;
  signal gl_ram_n_213, gl_ram_n_214, gl_ram_n_215, gl_ram_n_216, gl_ram_n_217 : std_logic;
  signal gl_ram_n_218, gl_ram_n_219, gl_ram_n_220, gl_ram_n_221, gl_ram_n_222 : std_logic;
  signal gl_ram_n_223, gl_ram_n_224, gl_ram_n_225, gl_ram_n_226, gl_ram_n_227 : std_logic;
  signal gl_ram_n_228, gl_ram_n_229, gl_ram_n_230, gl_ram_n_231, gl_ram_n_232 : std_logic;
  signal gl_ram_n_233, gl_ram_n_234, gl_ram_n_235, gl_ram_n_236, gl_ram_n_237 : std_logic;
  signal gl_ram_n_238, gl_ram_n_239, gl_ram_n_240, gl_ram_n_241, gl_ram_n_242 : std_logic;
  signal gl_ram_n_243, gl_ram_n_244, gl_ram_n_245, gl_ram_n_246, gl_ram_n_247 : std_logic;
  signal gl_ram_n_248, gl_ram_n_249, gl_ram_n_250, gl_ram_n_251, gl_ram_n_252 : std_logic;
  signal gl_ram_n_253, gl_ram_n_254, gl_ram_n_255, gl_ram_n_256, gl_ram_n_257 : std_logic;
  signal gl_ram_n_258, gl_ram_n_259, gl_ram_n_260, gl_ram_n_261, gl_ram_n_262 : std_logic;
  signal gl_ram_n_263, gl_ram_n_264, gl_ram_n_265, gl_ram_n_266, gl_ram_n_267 : std_logic;
  signal gl_ram_n_268, gl_ram_n_269, gl_ram_n_270, gl_ram_n_271, gl_ram_n_272 : std_logic;
  signal gl_ram_n_273, gl_ram_n_274, gl_ram_n_275, gl_ram_n_276, gl_ram_n_277 : std_logic;
  signal gl_ram_n_278, gl_ram_n_279, gl_ram_n_280, gl_ram_n_281, gl_ram_n_282 : std_logic;
  signal gl_ram_n_283, gl_ram_n_284, gl_ram_n_285, gl_ram_n_286, gl_ram_n_287 : std_logic;
  signal gl_ram_n_288, gl_ram_n_289, gl_ram_n_290, gl_ram_n_291, gl_ram_n_292 : std_logic;
  signal gl_ram_n_293, gl_ram_n_294, gl_ram_n_295, gl_ram_n_296, gl_ram_n_297 : std_logic;
  signal gl_ram_n_298, gl_ram_n_299, gl_ram_n_300, gl_ram_n_301, gl_ram_n_302 : std_logic;
  signal gl_ram_n_303, gl_ram_n_304, gl_ram_n_305, gl_ram_n_306, gl_ram_n_307 : std_logic;
  signal gl_ram_n_308, gl_ram_n_309, gl_ram_n_310, gl_ram_n_311, gl_ram_n_312 : std_logic;
  signal gl_ram_n_313, gl_ram_n_314, gl_ram_n_315, gl_ram_n_316, gl_ram_n_317 : std_logic;
  signal gl_ram_n_318, gl_ram_n_319, gl_ram_n_320, gl_ram_n_321, gl_ram_n_322 : std_logic;
  signal gl_ram_n_323, gl_ram_n_324, gl_ram_n_325, gl_ram_n_326, gl_ram_n_327 : std_logic;
  signal gl_ram_n_328, gl_ram_n_329, gl_ram_n_330, gl_ram_n_331, gl_ram_n_332 : std_logic;
  signal gl_ram_n_333, gl_ram_n_334, gl_ram_n_335, gl_ram_n_336, gl_ram_n_337 : std_logic;
  signal gl_ram_n_338, gl_ram_n_339, gl_ram_n_340, gl_ram_n_341, gl_ram_n_342 : std_logic;
  signal gl_ram_n_343, gl_ram_n_344, gl_ram_n_345, gl_ram_n_346, gl_ram_n_347 : std_logic;
  signal gl_ram_n_348, gl_ram_n_349, gl_ram_n_350, gl_ram_n_351, gl_ram_n_352 : std_logic;
  signal gl_ram_n_353, gl_ram_n_354, gl_ram_n_355, gl_ram_n_356, gl_ram_n_357 : std_logic;
  signal gl_ram_n_358, gl_ram_n_359, gl_ram_n_360, gl_ram_n_361, gl_ram_n_362 : std_logic;
  signal gl_ram_n_363, gl_ram_n_364, gl_ram_n_365, gl_ram_n_366, gl_ram_n_367 : std_logic;
  signal gl_ram_n_368, gl_ram_n_369, gl_ram_n_370, gl_ram_n_371, gl_ram_n_372 : std_logic;
  signal gl_ram_n_373, gl_ram_n_374, gl_ram_n_375, gl_ram_n_376, gl_ram_n_377 : std_logic;
  signal gl_ram_n_378, gl_ram_n_379, gl_ram_n_380, gl_ram_n_381, gl_ram_n_382 : std_logic;
  signal gl_ram_n_383, gl_ram_n_384, gl_ram_n_385, gl_ram_n_386, gl_ram_n_387 : std_logic;
  signal gl_ram_n_388, gl_ram_n_389, gl_ram_n_390, gl_ram_n_391, gl_ram_n_392 : std_logic;
  signal gl_ram_n_393, gl_ram_n_394, gl_ram_n_395, gl_ram_n_396, gl_ram_n_397 : std_logic;
  signal gl_ram_n_398, gl_ram_n_399, gl_ram_n_400, gl_ram_n_401, gl_ram_n_402 : std_logic;
  signal gl_ram_n_403, gl_ram_n_404, gl_ram_n_405, gl_ram_n_406, gl_ram_n_407 : std_logic;
  signal gl_ram_n_408, gl_ram_n_409, gl_ram_n_410, gl_ram_n_411, gl_ram_n_412 : std_logic;
  signal gl_ram_n_413, gl_ram_n_414, gl_ram_n_415, gl_ram_n_416, gl_ram_n_417 : std_logic;
  signal gl_ram_n_418, gl_ram_n_419, gl_ram_n_420, gl_ram_n_421, gl_ram_n_422 : std_logic;
  signal gl_ram_n_423, gl_ram_n_424, gl_ram_n_425, gl_ram_n_426, gl_ram_n_427 : std_logic;
  signal gl_ram_n_428, gl_ram_n_429, gl_ram_n_430, gl_ram_n_431, gl_ram_n_432 : std_logic;
  signal gl_ram_n_433, gl_ram_n_434, gl_ram_n_435, gl_ram_n_436, gl_ram_n_437 : std_logic;
  signal gl_ram_n_438, gl_ram_n_439, gl_ram_n_440, gl_ram_n_441, gl_ram_n_442 : std_logic;
  signal gl_ram_n_443, gl_ram_n_444, gl_ram_n_445, gl_ram_n_446, gl_ram_n_447 : std_logic;
  signal gl_ram_n_448, gl_ram_n_449, gl_ram_n_450, gl_ram_n_451, gl_ram_n_452 : std_logic;
  signal gl_ram_n_453, gl_ram_n_454, gl_ram_n_455, gl_ram_n_456, gl_ram_n_457 : std_logic;
  signal gl_ram_n_458, gl_ram_n_459, gl_ram_n_460, gl_ram_n_461, gl_ram_n_462 : std_logic;
  signal gl_ram_n_463, gl_ram_n_464, gl_ram_n_465, gl_ram_n_466, gl_ram_n_467 : std_logic;
  signal gl_ram_n_468, gl_ram_n_469, gl_ram_n_470, gl_ram_n_471, gl_ram_n_472 : std_logic;
  signal gl_ram_n_473, gl_ram_n_474, gl_ram_n_475, gl_ram_n_476, gl_ram_n_477 : std_logic;
  signal gl_ram_n_478, gl_ram_n_479, gl_ram_n_480, gl_ram_n_481, gl_ram_n_482 : std_logic;
  signal gl_ram_n_483, gl_ram_n_484, gl_ram_n_485, gl_ram_n_486, gl_ram_n_487 : std_logic;
  signal gl_ram_n_488, gl_ram_n_489, gl_ram_n_490, gl_ram_n_491, gl_ram_n_492 : std_logic;
  signal gl_ram_n_493, gl_ram_n_494, gl_ram_n_495, gl_ram_n_496, gl_ram_n_497 : std_logic;
  signal gl_ram_n_498, gl_ram_n_499, gl_ram_n_500, gl_ram_n_501, gl_ram_n_502 : std_logic;
  signal gl_ram_n_503, gl_ram_n_504, gl_ram_n_505, gl_ram_n_506, gl_ram_n_507 : std_logic;
  signal gl_ram_n_508, gl_ram_n_509, gl_ram_n_510, gl_ram_n_511, gl_ram_n_512 : std_logic;
  signal gl_ram_n_513, gl_ram_n_514, gl_ram_n_515, gl_ram_n_516, gl_ram_n_517 : std_logic;
  signal gl_ram_n_518, gl_ram_n_519, gl_ram_n_520, gl_ram_n_521, gl_ram_n_522 : std_logic;
  signal gl_ram_n_523, gl_ram_n_524, gl_ram_n_525, gl_ram_n_526, gl_ram_n_527 : std_logic;
  signal gl_ram_n_528, gl_ram_n_529, gl_ram_n_530, gl_ram_n_531, gl_ram_n_532 : std_logic;
  signal gl_ram_n_533, gl_ram_n_534, gl_ram_n_535, gl_ram_n_536, gl_ram_n_537 : std_logic;
  signal gl_ram_n_538, gl_ram_n_539, gl_ram_n_540, gl_ram_n_541, gl_ram_n_542 : std_logic;
  signal gl_ram_n_543, gl_ram_n_544, gl_ram_n_545, gl_ram_n_546, gl_ram_n_547 : std_logic;
  signal gl_ram_n_548, gl_ram_n_549, gl_ram_n_550, gl_ram_n_551, gl_ram_n_552 : std_logic;
  signal gl_ram_n_553, gl_ram_n_554, gl_ram_n_555, gl_ram_n_556, gl_ram_n_557 : std_logic;
  signal gl_ram_n_558, gl_ram_n_559, gl_ram_n_560, gl_ram_n_561, gl_ram_n_562 : std_logic;
  signal gl_ram_n_563, gl_ram_n_564, gl_ram_n_565, gl_ram_n_566, gl_ram_n_567 : std_logic;
  signal gl_ram_n_568, gl_ram_n_569, gl_ram_n_570, gl_ram_n_571, gl_ram_n_572 : std_logic;
  signal gl_ram_n_573, gl_ram_n_574, gl_ram_n_575, gl_ram_n_576, gl_ram_n_577 : std_logic;
  signal gl_ram_n_578, gl_ram_n_579, gl_ram_n_580, gl_ram_n_581, gl_ram_n_582 : std_logic;
  signal gl_ram_n_583, gl_ram_n_584, gl_ram_n_585, gl_ram_n_586, gl_ram_n_587 : std_logic;
  signal gl_ram_n_588, gl_ram_n_589, gl_ram_n_590, gl_ram_n_591, gl_ram_n_592 : std_logic;
  signal gl_ram_n_593, gl_ram_n_594, gl_ram_n_595, gl_ram_n_596, gl_ram_n_597 : std_logic;
  signal gl_ram_n_598, gl_ram_n_599, gl_ram_n_600, gl_ram_n_601, gl_ram_n_602 : std_logic;
  signal gl_ram_n_603, gl_ram_n_604, gl_ram_n_605, gl_ram_n_606, gl_ram_n_607 : std_logic;
  signal gl_ram_n_608, gl_ram_n_609, gl_ram_n_610, gl_ram_n_611, gl_ram_n_612 : std_logic;
  signal gl_ram_n_613, gl_ram_n_614, gl_ram_n_615, gl_ram_n_616, gl_ram_n_617 : std_logic;
  signal gl_ram_n_618, gl_ram_n_619, gl_ram_n_620, gl_ram_n_621, gl_ram_n_622 : std_logic;
  signal gl_ram_n_623, gl_ram_n_624, gl_ram_n_625, gl_ram_n_626, gl_ram_n_627 : std_logic;
  signal gl_ram_n_628, gl_ram_n_629, gl_ram_n_630, gl_ram_n_631, gl_ram_n_632 : std_logic;
  signal gl_ram_n_633, gl_ram_n_634, gl_ram_n_635, gl_ram_n_636, gl_ram_n_637 : std_logic;
  signal gl_ram_n_638, gl_ram_n_639, gl_ram_n_640, gl_ram_n_641, gl_ram_n_642 : std_logic;
  signal gl_ram_n_643, gl_ram_n_644, gl_ram_n_645, gl_ram_n_646, gl_ram_n_647 : std_logic;
  signal gl_ram_n_648, gl_ram_n_649, gl_ram_n_650, gl_ram_n_651, gl_ram_n_652 : std_logic;
  signal gl_ram_n_653, gl_ram_n_654, gl_ram_n_655, gl_ram_n_656, gl_ram_n_657 : std_logic;
  signal gl_ram_n_658, gl_ram_n_659, gl_ram_n_660, gl_ram_n_661, gl_ram_n_662 : std_logic;
  signal gl_ram_n_663, gl_ram_n_664, gl_ram_n_665, gl_ram_n_666, gl_ram_n_667 : std_logic;
  signal gl_ram_n_668, gl_ram_n_669, gl_ram_n_670, gl_ram_n_671, gl_ram_n_672 : std_logic;
  signal gl_ram_n_673, gl_ram_n_674, gl_ram_n_675, gl_ram_n_676, gl_ram_n_677 : std_logic;
  signal gl_ram_n_678, gl_ram_n_679, gl_ram_n_680, gl_ram_n_681, gl_ram_n_682 : std_logic;
  signal gl_ram_n_683, gl_ram_n_684, gl_ram_n_685, gl_ram_n_686, gl_ram_n_687 : std_logic;
  signal gl_ram_n_688, gl_ram_n_689, gl_ram_n_690, gl_ram_n_691, gl_ram_n_692 : std_logic;
  signal gl_ram_n_693, gl_ram_n_694, gl_ram_n_695, gl_ram_n_696, gl_ram_n_697 : std_logic;
  signal gl_ram_n_698, gl_ram_n_699, gl_ram_n_700, gl_ram_n_701, gl_ram_n_702 : std_logic;
  signal gl_ram_n_703, gl_ram_n_704, gl_ram_n_705, gl_ram_n_706, gl_ram_n_707 : std_logic;
  signal gl_ram_n_708, gl_ram_n_709, gl_ram_n_710, gl_ram_n_711, gl_ram_n_712 : std_logic;
  signal gl_ram_n_713, gl_ram_n_714, gl_ram_n_715, gl_ram_n_716, gl_ram_n_717 : std_logic;
  signal gl_ram_n_718, gl_ram_n_719, gl_ram_n_720, gl_ram_n_721, gl_ram_n_722 : std_logic;
  signal gl_ram_n_723, gl_ram_n_724, gl_ram_n_725, gl_ram_n_726, gl_ram_n_727 : std_logic;
  signal gl_ram_n_728, gl_ram_n_729, gl_ram_n_730, gl_ram_n_731, gl_ram_n_732 : std_logic;
  signal gl_ram_n_733, gl_ram_n_734, gl_ram_n_735, gl_ram_n_736, gl_ram_n_737 : std_logic;
  signal gl_ram_n_738, gl_ram_n_739, gl_ram_n_740, gl_ram_n_741, gl_ram_n_742 : std_logic;
  signal gl_ram_n_743, gl_ram_n_744, gl_ram_n_745, gl_ram_n_746, gl_ram_n_747 : std_logic;
  signal gl_ram_n_748, gl_ram_n_749, gl_ram_n_750, gl_ram_n_751, gl_ram_n_752 : std_logic;
  signal gl_ram_n_753, gl_ram_n_754, gl_ram_n_755, gl_ram_n_756, gl_ram_n_757 : std_logic;
  signal gl_ram_n_758, gl_ram_n_759, gl_ram_n_760, gl_ram_n_761, gl_ram_n_762 : std_logic;
  signal gl_ram_n_763, gl_ram_n_764, gl_ram_n_765, gl_ram_n_766, gl_ram_n_767 : std_logic;
  signal gl_ram_n_768, gl_ram_n_769, gl_ram_n_770, gl_ram_n_771, gl_ram_n_772 : std_logic;
  signal gl_ram_n_773, gl_ram_n_774, gl_ram_n_775, gl_ram_n_776, gl_ram_n_777 : std_logic;
  signal gl_ram_n_778, gl_ram_n_779, gl_ram_n_780, gl_ram_n_781, gl_ram_n_782 : std_logic;
  signal gl_ram_n_783, gl_ram_n_784, gl_ram_n_785, gl_ram_n_786, gl_ram_n_787 : std_logic;
  signal gl_ram_n_788, gl_ram_n_789, gl_ram_n_790, gl_ram_n_791, gl_ram_n_792 : std_logic;
  signal gl_ram_n_793, gl_ram_n_794, gl_ram_n_795, gl_ram_n_796, gl_ram_n_797 : std_logic;
  signal gl_ram_n_798, gl_ram_n_799, gl_ram_n_800, gl_ram_n_801, gl_ram_n_802 : std_logic;
  signal gl_ram_n_803, gl_ram_n_804, gl_ram_n_805, gl_ram_n_806, gl_ram_n_807 : std_logic;
  signal gl_ram_n_808, gl_ram_n_809, gl_ram_n_810, gl_ram_n_811, gl_ram_n_812 : std_logic;
  signal gl_ram_n_813, gl_ram_n_814, gl_ram_n_815, gl_ram_n_816, gl_ram_n_817 : std_logic;
  signal gl_ram_n_818, gl_ram_n_819, gl_ram_n_820, gl_ram_n_821, gl_ram_n_822 : std_logic;
  signal gl_ram_n_823, gl_ram_n_824, gl_ram_n_825, gl_ram_n_826, gl_rom_n_0 : std_logic;
  signal gl_rom_n_1, gl_rom_n_2, gl_rom_n_3, gl_rom_n_4, gl_rom_n_5 : std_logic;
  signal gl_rom_n_6, gl_rom_n_7, gl_rom_n_8, gl_rom_n_9, gl_rom_n_10 : std_logic;
  signal gl_rom_n_11, gl_rom_n_12, gl_rom_n_13, gl_rom_n_14, gl_rom_n_15 : std_logic;
  signal gl_rom_n_16, gl_rom_n_17, gl_rom_n_18, gl_rom_n_19, gl_rom_n_20 : std_logic;
  signal gl_rom_n_21, gl_rom_n_22, gl_rom_n_23, gl_rom_n_24, gl_rom_n_25 : std_logic;
  signal gl_rom_n_26, gl_rom_n_27, gl_rom_n_28, gl_rom_n_29, gl_rom_n_30 : std_logic;
  signal gl_rom_n_31, gl_rom_n_32, gl_rom_n_33, gl_rom_n_34, gl_rom_n_35 : std_logic;
  signal gl_rom_n_36, gl_rom_n_37, gl_rom_n_38, gl_rom_n_39, gl_rom_n_40 : std_logic;
  signal gl_rom_n_41, gl_rom_n_42, gl_rom_n_43, gl_rom_n_44, gl_rom_n_45 : std_logic;
  signal gl_rom_n_46, gl_rom_n_47, gl_rom_n_48, gl_rom_n_49, gl_rom_n_50 : std_logic;
  signal gl_rom_n_51, gl_rom_n_52, gl_rom_n_53, gl_rom_n_54, gl_rom_n_55 : std_logic;
  signal gl_rom_n_56, gl_rom_n_57, gl_rom_n_58, gl_rom_n_59, gl_rom_n_60 : std_logic;
  signal gl_rom_n_61, gl_rom_n_62, gl_rom_n_63, gl_rom_n_64, gl_rom_n_65 : std_logic;
  signal gl_rom_n_66, gl_rom_n_67, gl_rom_n_68, gl_rom_n_69, gl_rom_n_70 : std_logic;
  signal gl_rom_n_71, gl_rom_n_72, gl_rom_n_73, gl_rom_n_74, gl_rom_n_75 : std_logic;
  signal gl_rom_n_76, gl_rom_n_77, gl_rom_n_78, gl_rom_n_79, gl_rom_n_80 : std_logic;
  signal gl_rom_n_81, gl_rom_n_82, gl_rom_n_83, gl_rom_n_84, gl_rom_n_85 : std_logic;
  signal gl_rom_n_86, gl_rom_n_87, gl_rom_n_88, gl_rom_n_89, gl_rom_n_90 : std_logic;
  signal gl_rom_n_91, gl_rom_n_92, gl_rom_n_93, gl_rom_n_94, gl_rom_n_95 : std_logic;
  signal gl_rom_n_96, gl_rom_n_97, gl_rom_n_98, gl_rom_n_99, gl_rom_n_100 : std_logic;
  signal gl_rom_n_101, gl_rom_n_102, gl_rom_n_103, gl_rom_n_104, gl_rom_n_105 : std_logic;
  signal gl_rom_n_106, gl_rom_n_107, gl_rom_n_108, gl_rom_n_109, gl_rom_n_110 : std_logic;
  signal gl_rom_n_111, gl_rom_n_112, gl_rom_n_113, gl_rom_n_114, gl_rom_n_115 : std_logic;
  signal gl_rom_n_116, gl_rom_n_117, gl_rom_n_118, gl_rom_n_119, gl_rom_n_120 : std_logic;
  signal gl_rom_n_121, gl_rom_n_122, gl_rom_n_123, gl_rom_n_124, gl_rom_n_125 : std_logic;
  signal gl_rom_n_126, gl_rom_n_127, gl_rom_n_128, gl_rom_n_129, gl_rom_n_130 : std_logic;
  signal gl_rom_n_131, gl_rom_n_132, gl_rom_n_133, gl_rom_n_134, gl_rom_n_135 : std_logic;
  signal gl_rom_n_136, gl_rom_n_137, gl_rom_n_138, gl_rom_n_139, gl_rom_n_140 : std_logic;
  signal gl_rom_n_141, gl_rom_n_142, gl_rom_n_143, gl_rom_n_144, gl_rom_n_145 : std_logic;
  signal gl_rom_n_146, gl_rom_n_147, gl_rom_n_148, gl_rom_n_149, gl_rom_n_150 : std_logic;
  signal gl_rom_n_151, gl_rom_n_152, gl_rom_n_153, gl_rom_n_154, gl_rom_n_155 : std_logic;
  signal gl_rom_n_156, gl_rom_n_157, gl_rom_n_158, gl_rom_n_159, gl_rom_n_160 : std_logic;
  signal gl_rom_n_161, gl_rom_n_162, gl_rom_n_163, gl_rom_n_164, gl_rom_n_165 : std_logic;
  signal gl_rom_n_166, gl_rom_n_167, gl_rom_n_168, gl_rom_n_169, gl_rom_n_170 : std_logic;
  signal gl_rom_n_171, gl_rom_n_172, gl_rom_n_173, gl_rom_n_174, gl_rom_n_175 : std_logic;
  signal gl_rom_n_176, gl_rom_n_177, gl_rom_n_178, gl_rom_n_179, gl_rom_n_180 : std_logic;
  signal gl_rom_n_181, gl_rom_n_182, gl_rom_n_183, gl_rom_n_184, gl_rom_n_185 : std_logic;
  signal gl_rom_n_186, gl_rom_n_187, gl_rom_n_188, gl_rom_n_189, gl_rom_n_190 : std_logic;
  signal gl_rom_n_191, gl_rom_n_192, gl_rom_n_193, gl_rom_n_194, gl_rom_n_195 : std_logic;
  signal gl_rom_n_196, gl_rom_n_197, gl_rom_n_198, gl_rom_n_199, gl_rom_n_200 : std_logic;
  signal gl_rom_n_201, gl_rom_n_202, gl_rom_n_203, gl_rom_n_204, gl_rom_n_205 : std_logic;
  signal gl_rom_n_206, gl_rom_n_207, gl_rom_n_208, gl_rom_n_209, gl_rom_n_210 : std_logic;
  signal gl_rom_n_211, gl_rom_n_212, gl_rom_n_213, gl_rom_n_214, gl_rom_n_215 : std_logic;
  signal gl_rom_n_216, gl_rom_n_217, gl_rom_n_218, gl_rom_n_219, gl_rom_n_220 : std_logic;
  signal gl_rom_n_221, gl_rom_n_222, gl_rom_n_223, gl_rom_n_224, gl_rom_n_225 : std_logic;
  signal gl_rom_n_226, gl_rom_n_227, gl_rom_n_228, gl_rom_n_229, gl_rom_n_230 : std_logic;
  signal gl_rom_n_231, gl_rom_n_232, gl_rom_n_233, gl_rom_n_234, gl_rom_n_235 : std_logic;
  signal gl_rom_n_236, gl_rom_n_237, gl_rom_n_238, gl_rom_n_239, gl_rom_n_240 : std_logic;
  signal gl_rom_n_241, gl_rom_n_242, gl_rom_n_243, gl_rom_n_244, gl_rom_n_245 : std_logic;
  signal gl_rom_n_246, gl_rom_n_247, gl_rom_n_248, gl_rom_n_249, gl_rom_n_250 : std_logic;
  signal gl_rom_n_251, gl_rom_n_252, gl_rom_n_253, gl_rom_n_254, gl_rom_n_255 : std_logic;
  signal gl_rom_n_256, gl_rom_n_257, gl_rom_n_258, gl_rom_n_259, gl_rom_n_260 : std_logic;
  signal gl_rom_n_261, gl_rom_n_262, gl_rom_n_263, gl_rom_n_264, gl_rom_n_265 : std_logic;
  signal gl_rom_n_266, gl_rom_n_267, gl_rom_n_268, gl_rom_n_269, gl_rom_n_270 : std_logic;
  signal gl_rom_n_271, gl_rom_n_272, gl_rom_n_273, gl_rom_n_274, gl_rom_n_275 : std_logic;
  signal gl_rom_n_276, gl_rom_n_277, gl_rom_n_278, gl_rom_n_279, gl_rom_n_280 : std_logic;
  signal gl_rom_n_281, gl_rom_n_282, gl_rom_n_283, gl_rom_n_284, gl_rom_n_285 : std_logic;
  signal gl_rom_n_286, gl_rom_n_287, gl_rom_n_288, gl_rom_n_289, gl_rom_n_290 : std_logic;
  signal gl_rom_n_291, gl_rom_n_292, gl_rom_n_293, gl_rom_n_294, gl_rom_n_295 : std_logic;
  signal gl_rom_n_296, gl_rom_n_297, gl_rom_n_298, gl_rom_n_299, gl_rom_n_300 : std_logic;
  signal gl_rom_n_301, gl_rom_n_302, gl_rom_n_303, gl_rom_n_304, gl_rom_n_305 : std_logic;
  signal gl_rom_n_306, gl_rom_n_307, gl_rom_n_308, gl_rom_n_309, gl_rom_n_310 : std_logic;
  signal gl_rom_n_311, gl_rom_n_312, gl_rom_n_313, gl_rom_n_314, gl_rom_n_315 : std_logic;
  signal gl_rom_n_316, gl_rom_n_317, gl_rom_n_318, gl_rom_n_319, gl_rom_n_320 : std_logic;
  signal gl_rom_n_321, gl_rom_n_322, gl_rom_n_323, gl_rom_n_324, gl_rom_n_325 : std_logic;
  signal gl_rom_n_326, gl_rom_n_327, gl_rom_n_328, gl_rom_n_329, gl_rom_n_330 : std_logic;
  signal gl_rom_n_331, gl_rom_n_332, gl_rom_n_333, gl_rom_n_334, gl_rom_n_335 : std_logic;
  signal gl_rom_n_336, gl_rom_n_337, gl_rom_n_338, gl_rom_n_339, gl_rom_n_340 : std_logic;
  signal gl_rom_n_341, gl_rom_n_342, gl_rom_n_343, gl_rom_n_344, gl_rom_n_345 : std_logic;
  signal gl_rom_n_346, gl_rom_n_347, gl_rom_n_348, gl_rom_n_349, gl_rom_n_350 : std_logic;
  signal gl_rom_n_351, gl_rom_n_352, gl_rom_n_353, gl_rom_n_354, gl_rom_n_355 : std_logic;
  signal gl_rom_n_356, gl_rom_n_357, gl_rom_n_358, gl_rom_n_359, gl_rom_n_360 : std_logic;
  signal gl_rom_n_361, gl_rom_n_362, gl_rom_n_363, gl_rom_n_364, gl_rom_n_365 : std_logic;
  signal gl_rom_n_366, gl_rom_n_367, gl_rom_n_368, gl_rom_n_369, gl_rom_n_370 : std_logic;
  signal gl_rom_n_371, gl_rom_n_372, gl_rom_n_373, gl_rom_n_374, gl_rom_n_375 : std_logic;
  signal gl_rom_n_376, gl_rom_n_377, gl_rom_n_378, gl_rom_n_379, gl_rom_n_380 : std_logic;
  signal gl_rom_n_381, gl_rom_n_382, gl_rom_n_383, gl_rom_n_384, gl_rom_n_385 : std_logic;
  signal gl_rom_n_386, gl_rom_n_387, gl_rom_n_388, gl_rom_n_389, gl_rom_n_390 : std_logic;
  signal gl_rom_n_391, gl_rom_n_392, gl_rom_n_393, gl_rom_n_394, gl_rom_n_395 : std_logic;
  signal gl_rom_n_396, gl_rom_n_397, gl_rom_n_398, gl_rom_n_399, gl_rom_n_400 : std_logic;
  signal gl_rom_n_401, gl_rom_n_402, gl_rom_n_403, gl_rom_n_404, gl_rom_n_405 : std_logic;
  signal gl_rom_n_406, gl_rom_n_407, gl_rom_n_408, gl_rom_n_409, gl_rom_n_410 : std_logic;
  signal gl_rom_n_411, gl_rom_n_412, gl_rom_n_413, gl_rom_n_414, gl_rom_n_415 : std_logic;
  signal gl_rom_n_416, gl_rom_n_417, gl_rom_n_418, gl_rom_n_419, gl_rom_n_420 : std_logic;
  signal gl_rom_n_421, gl_rom_n_422, gl_rom_n_423, gl_rom_n_424, gl_rom_n_425 : std_logic;
  signal gl_rom_n_426, gl_rom_n_427, gl_rom_n_428, gl_rom_n_429, gl_rom_n_430 : std_logic;
  signal gl_rom_n_431, gl_rom_n_432, gl_rom_n_433, gl_rom_n_434, gl_rom_n_435 : std_logic;
  signal gl_rom_n_436, gl_rom_n_437, gl_rom_n_438, gl_rom_n_439, gl_rom_n_440 : std_logic;
  signal gl_rom_n_441, gl_rom_n_442, gl_rom_n_443, gl_rom_n_444, gl_rom_n_445 : std_logic;
  signal gl_rom_n_446, gl_rom_n_447, gl_rom_n_448, gl_rom_n_449, gl_rom_n_450 : std_logic;
  signal gl_rom_n_451, gl_rom_n_452, gl_rom_n_453, gl_rom_n_454, gl_rom_n_455 : std_logic;
  signal gl_rom_n_456, gl_rom_n_457, gl_rom_n_458, gl_rom_n_459, gl_rom_n_460 : std_logic;
  signal gl_rom_n_461, gl_rom_n_462, gl_rom_n_463, gl_rom_n_464, gl_rom_n_465 : std_logic;
  signal gl_rom_n_466, gl_rom_n_467, gl_rom_n_468, gl_rom_n_469, gl_rom_n_470 : std_logic;
  signal gl_rom_n_471, gl_rom_n_472, gl_rom_n_473, gl_rom_n_474, gl_rom_n_475 : std_logic;
  signal gl_rom_n_476, gl_rom_n_477, gl_rom_n_478, gl_rom_n_479, gl_rom_n_480 : std_logic;
  signal gl_rom_n_481, gl_rom_n_482, gl_rom_n_483, gl_rom_n_484, gl_rom_n_485 : std_logic;
  signal gl_rom_n_486, gl_rom_n_487, gl_rom_n_488, gl_rom_n_489, gl_rom_n_490 : std_logic;
  signal gl_rom_n_491, gl_rom_n_492, gl_rom_n_493, gl_rom_n_494, gl_rom_n_495 : std_logic;
  signal gl_rom_n_496, gl_rom_n_497, gl_rom_n_498, gl_rom_n_499, gl_rom_n_500 : std_logic;
  signal gl_rom_n_501, gl_rom_n_502, gl_rom_n_503, gl_rom_n_504, gl_rom_n_505 : std_logic;
  signal gl_rom_n_506, gl_rom_n_507, gl_rom_n_508, gl_rom_n_509, gl_rom_n_510 : std_logic;
  signal gl_rom_n_511, gl_rom_n_512, gl_rom_n_513, gl_rom_n_514, gl_rom_n_515 : std_logic;
  signal gl_rom_n_516, gl_rom_n_517, gl_rom_n_518, gl_rom_n_519, gl_rom_n_520 : std_logic;
  signal gl_rom_n_521, gl_rom_n_522, gl_rom_n_523, gl_rom_n_524, gl_rom_n_525 : std_logic;
  signal gl_rom_n_526, gl_rom_n_527, gl_rom_n_528, gl_rom_n_529, gl_rom_n_530 : std_logic;
  signal gl_rom_n_531, gl_rom_n_532, gl_rom_n_533, gl_rom_n_534, gl_rom_n_535 : std_logic;
  signal gl_rom_n_536, gl_rom_n_537, gl_rom_n_538, gl_rom_n_539, gl_rom_n_540 : std_logic;
  signal gl_rom_n_541, gl_rom_n_542, gl_rom_n_543, gl_rom_n_544, gl_rom_n_545 : std_logic;
  signal gl_rom_n_546, gl_rom_n_547, gl_rom_n_548, gl_rom_n_549, gl_rom_n_550 : std_logic;
  signal gl_rom_n_551, gl_rom_n_552, gl_rom_n_553, gl_rom_n_554, gl_rom_n_555 : std_logic;
  signal gl_rom_n_556, gl_rom_n_557, gl_rom_n_558, gl_rom_n_559, gl_rom_n_560 : std_logic;
  signal gl_rom_n_561, gl_rom_n_562, gl_rom_n_563, gl_rom_n_564, gl_rom_n_565 : std_logic;
  signal gl_rom_n_566, gl_rom_n_567, gl_rom_n_568, gl_rom_n_569, gl_rom_n_570 : std_logic;
  signal gl_rom_n_571, gl_rom_n_572, gl_rom_n_573, gl_rom_n_574, gl_rom_n_575 : std_logic;
  signal gl_rom_n_576, gl_rom_n_577, gl_rom_n_578, gl_rom_n_579, gl_rom_n_580 : std_logic;
  signal gl_rom_n_581, gl_rom_n_582, gl_rom_n_583, gl_rom_n_584, gl_rom_n_585 : std_logic;
  signal gl_rom_n_586, gl_rom_n_587, gl_rom_n_588, gl_rom_n_589, gl_rom_n_590 : std_logic;
  signal gl_rom_n_591, gl_rom_n_592, gl_rom_n_593, gl_rom_n_594, gl_rom_n_595 : std_logic;
  signal gl_rom_n_596, gl_rom_n_597, gl_rom_n_598, gl_rom_n_599, gl_rom_n_600 : std_logic;
  signal gl_rom_n_601, gl_rom_n_602, gl_rom_n_603, gl_rom_n_604, gl_rom_n_605 : std_logic;
  signal gl_rom_n_606, gl_rom_n_607, gl_rom_n_608, gl_rom_n_609, gl_rom_n_610 : std_logic;
  signal gl_rom_n_611, gl_rom_n_612, gl_rom_n_613, gl_rom_n_614, gl_rom_n_615 : std_logic;
  signal gl_rom_n_616, gl_rom_n_617, gl_rom_n_618, gl_rom_n_619, gl_rom_n_620 : std_logic;
  signal gl_rom_n_621, gl_rom_n_622, gl_rom_n_623, gl_rom_n_624, gl_rom_n_625 : std_logic;
  signal gl_rom_n_626, gl_rom_n_627, gl_rom_n_628, gl_rom_n_629, gl_rom_n_630 : std_logic;
  signal gl_rom_n_631, gl_rom_n_632, gl_rom_n_633, gl_rom_n_634, gl_rom_n_635 : std_logic;
  signal gl_rom_n_636, gl_rom_n_637, gl_rom_n_638, gl_rom_n_639, gl_rom_n_640 : std_logic;
  signal gl_rom_n_641, gl_rom_n_642, gl_rom_n_643, gl_rom_n_644, gl_rom_n_645 : std_logic;
  signal gl_rom_n_646, gl_rom_n_647, gl_rom_n_648, gl_rom_n_649, gl_rom_n_650 : std_logic;
  signal gl_rom_n_651, gl_rom_n_652, gl_rom_n_653, gl_rom_n_654, gl_rom_n_655 : std_logic;
  signal gl_rom_n_656, gl_rom_n_657, gl_rom_n_658, gl_rom_n_659, gl_rom_n_660 : std_logic;
  signal gl_rom_n_661, gl_rom_n_662, gl_rom_n_663, gl_rom_n_664, gl_rom_n_665 : std_logic;
  signal gl_rom_n_666, gl_rom_n_667, gl_rom_n_668, gl_rom_n_669, gl_rom_n_670 : std_logic;
  signal gl_rom_n_671, gl_rom_n_672, gl_rom_n_673, gl_rom_n_674, gl_rom_n_675 : std_logic;
  signal gl_rom_n_676, gl_rom_n_677, gl_rom_n_678, gl_rom_n_679, gl_rom_n_680 : std_logic;
  signal gl_rom_n_681, gl_rom_n_682, gl_rom_n_683, gl_rom_n_684, gl_rom_n_685 : std_logic;
  signal gl_rom_n_686, gl_rom_n_687, gl_rom_n_688, gl_rom_n_689, gl_rom_n_690 : std_logic;
  signal gl_rom_n_691, gl_rom_n_692, gl_rom_n_693, gl_rom_n_694, gl_rom_n_695 : std_logic;
  signal gl_rom_n_696, gl_rom_n_697, gl_rom_n_698, gl_rom_n_699, gl_rom_n_700 : std_logic;
  signal gl_rom_n_701, gl_rom_n_702, gl_rom_n_703, gl_rom_n_704, gl_rom_n_705 : std_logic;
  signal gl_rom_n_706, gl_rom_n_707, gl_rom_n_708, gl_rom_n_709, gl_rom_n_710 : std_logic;
  signal gl_rom_n_711, gl_rom_n_712, gl_rom_n_713, gl_rom_n_714, gl_rom_n_715 : std_logic;
  signal gl_rom_n_716, gl_rom_n_717, gl_rom_n_718, gl_rom_n_719, gl_rom_n_720 : std_logic;
  signal gl_rom_n_721, gl_rom_n_722, gl_rom_n_723, gl_rom_n_724, gl_rom_n_725 : std_logic;
  signal gl_rom_n_726, gl_rom_n_727, gl_rom_n_728, gl_rom_n_729, gl_rom_n_730 : std_logic;
  signal gl_rom_n_731, gl_rom_n_732, gl_rom_n_733, gl_rom_n_734, gl_rom_n_735 : std_logic;
  signal gl_rom_n_736, gl_rom_n_737, gl_rom_n_738, gl_rom_n_739, gl_rom_n_740 : std_logic;
  signal gl_rom_n_741, gl_rom_n_742, gl_rom_n_743, gl_rom_n_744, gl_rom_n_745 : std_logic;
  signal gl_rom_n_746, gl_rom_n_747, gl_rom_n_748, gl_rom_n_749, gl_rom_n_750 : std_logic;
  signal gl_rom_n_751, gl_rom_n_752, gl_rom_n_753, gl_rom_n_754, gl_rom_n_755 : std_logic;
  signal gl_rom_n_756, gl_rom_n_757, gl_rom_n_758, gl_rom_n_759, gl_rom_n_760 : std_logic;
  signal gl_rom_n_761, gl_rom_n_762, gl_rom_n_763, gl_rom_n_764, gl_rom_n_765 : std_logic;
  signal gl_rom_n_766, gl_rom_n_767, gl_rom_n_768, gl_rom_n_769, gl_rom_n_770 : std_logic;
  signal gl_rom_n_771, gl_rom_n_772, gl_rom_n_773, gl_rom_n_774, gl_rom_n_775 : std_logic;
  signal gl_rom_n_776, gl_rom_n_777, gl_rom_n_778, gl_rom_n_779, gl_rom_n_780 : std_logic;
  signal gl_rom_n_781, gl_rom_n_782, gl_rom_n_783, gl_rom_n_784, gl_rom_n_785 : std_logic;
  signal gl_rom_n_786, gl_rom_n_787, gl_rom_n_788, gl_rom_n_789, gl_rom_n_790 : std_logic;
  signal gl_rom_n_791, gl_rom_n_792, gl_rom_n_793, gl_rom_n_794, gl_rom_n_795 : std_logic;
  signal gl_rom_n_796, gl_rom_n_797, gl_rom_n_798, gl_rom_n_799, gl_rom_n_800 : std_logic;
  signal gl_rom_n_801, gl_rom_n_802, gl_rom_n_803, gl_rom_n_804, gl_rom_n_805 : std_logic;
  signal gl_rom_n_806, gl_rom_n_807, gl_rom_n_808, gl_rom_n_809, gl_rom_n_810 : std_logic;
  signal gl_rom_n_811, gl_rom_n_812, gl_rom_n_813, gl_rom_n_814, gl_rom_n_815 : std_logic;
  signal gl_rom_n_816, gl_rom_n_817, gl_rom_n_818, gl_rom_n_819, gl_rom_n_820 : std_logic;
  signal gl_rom_n_821, gl_rom_n_822, gl_rom_n_823, gl_rom_n_824, gl_rom_n_825 : std_logic;
  signal gl_rom_n_826, gl_rom_n_827, gl_rom_n_828, gl_rom_n_829, gl_rom_n_830 : std_logic;
  signal gl_rom_n_831, gl_rom_n_832, gl_rom_n_833, gl_rom_n_834, gl_rom_n_835 : std_logic;
  signal gl_rom_n_836, gl_rom_n_837, gl_rom_n_838, gl_rom_n_839, gl_rom_n_840 : std_logic;
  signal gl_rom_n_841, gl_rom_n_842, gl_rom_n_843, gl_rom_n_844, gl_rom_n_845 : std_logic;
  signal gl_rom_n_846, gl_rom_n_847, gl_rom_n_848, gl_rom_n_849, gl_rom_n_850 : std_logic;
  signal gl_rom_n_851, gl_rom_n_852, gl_rom_n_853, gl_rom_n_854, gl_rom_n_855 : std_logic;
  signal gl_rom_n_856, gl_rom_n_857, gl_rom_n_858, gl_rom_n_859, gl_rom_n_860 : std_logic;
  signal gl_rom_n_861, gl_rom_n_862, gl_rom_n_863, gl_rom_n_864, gl_rom_n_865 : std_logic;
  signal gl_rom_n_866, gl_rom_n_867, gl_rom_n_868, gl_rom_n_869, gl_rom_n_870 : std_logic;
  signal gl_rom_n_871, gl_rom_n_872, gl_rom_n_873, gl_rom_n_874, gl_rom_n_875 : std_logic;
  signal gl_rom_n_876, gl_rom_n_877, gl_rom_n_878, gl_rom_n_879, gl_rom_n_880 : std_logic;
  signal gl_rom_n_881, gl_rom_n_882, gl_rom_n_883, gl_rom_n_884, gl_rom_n_885 : std_logic;
  signal gl_rom_n_886, gl_rom_n_887, gl_rom_n_888, gl_rom_n_889, gl_rom_n_890 : std_logic;
  signal gl_rom_n_891, gl_rom_n_892, gl_rom_n_893, gl_rom_n_894, gl_rom_n_895 : std_logic;
  signal gl_rom_n_896, gl_rom_n_897, gl_rom_n_898, gl_rom_n_899, gl_rom_n_900 : std_logic;
  signal gl_rom_n_901, gl_rom_n_902, gl_rom_n_903, gl_rom_n_904, gl_rom_n_905 : std_logic;
  signal gl_rom_n_906, gl_rom_n_907, gl_rom_n_908, gl_rom_n_909, gl_rom_n_910 : std_logic;
  signal gl_rom_n_911, gl_rom_n_912, gl_rom_n_913, gl_rom_n_914, gl_rom_n_915 : std_logic;
  signal gl_rom_n_916, gl_rom_n_917, gl_rom_n_918, gl_rom_n_919, gl_rom_n_920 : std_logic;
  signal gl_rom_n_921, gl_rom_n_922, gl_rom_n_923, gl_rom_n_924, gl_rom_n_925 : std_logic;
  signal gl_rom_n_926, gl_rom_n_927, gl_rom_n_928, gl_rom_n_929, gl_rom_n_930 : std_logic;
  signal gl_rom_n_931, gl_rom_n_932, gl_rom_n_933, gl_rom_n_934, gl_rom_n_935 : std_logic;
  signal gl_rom_n_936, gl_rom_n_937, gl_rom_n_938, gl_rom_n_939, gl_rom_n_940 : std_logic;
  signal gl_rom_n_941, gl_rom_n_942, gl_rom_n_943, gl_rom_n_944, gl_rom_n_945 : std_logic;
  signal gl_rom_n_946, gl_rom_n_947, gl_rom_n_948, gl_rom_n_949, gl_rom_n_950 : std_logic;
  signal gl_rom_n_951, gl_rom_n_952, gl_rom_n_953, gl_rom_n_954, gl_rom_n_955 : std_logic;
  signal gl_rom_n_956, gl_rom_n_957, gl_rom_n_958, gl_rom_n_959, gl_rom_n_960 : std_logic;
  signal gl_rom_n_961, gl_rom_n_962, gl_rom_n_963, gl_rom_n_964, gl_rom_n_965 : std_logic;
  signal gl_rom_n_966, gl_rom_n_967, gl_rom_n_968, gl_rom_n_969, gl_rom_n_970 : std_logic;
  signal gl_rom_n_971, gl_rom_n_972, gl_rom_n_973, gl_rom_n_974, gl_rom_n_975 : std_logic;
  signal gl_rom_n_976, gl_rom_n_977, gl_rom_n_978, gl_rom_n_979, gl_rom_n_980 : std_logic;
  signal gl_rom_n_981, gl_rom_n_982, gl_rom_n_983, gl_rom_n_984, gl_rom_n_985 : std_logic;
  signal gl_rom_n_986, gl_rom_n_987, gl_rom_n_988, gl_rom_n_989, gl_rom_n_990 : std_logic;
  signal gl_rom_n_991, gl_rom_n_992, gl_rom_n_993, gl_rom_n_994, gl_rom_n_995 : std_logic;
  signal gl_rom_n_996, gl_rom_n_997, gl_rom_n_998, gl_rom_n_999, gl_rom_n_1000 : std_logic;
  signal gl_rom_n_1001, gl_rom_n_1002, gl_rom_n_1003, gl_rom_n_1004, gl_rom_n_1005 : std_logic;
  signal gl_rom_n_1006, gl_rom_n_1007, gl_rom_n_1008, gl_rom_n_1009, gl_rom_n_1010 : std_logic;
  signal gl_rom_n_1011, gl_rom_n_1012, gl_rom_n_1013, gl_rom_n_1014, gl_rom_n_1015 : std_logic;
  signal gl_rom_n_1016, gl_rom_n_1017, gl_rom_n_1018, gl_rom_n_1019, gl_rom_n_1020 : std_logic;
  signal gl_rom_n_1021, gl_rom_n_1022, gl_rom_n_1023, gl_rom_n_1024, gl_rom_n_1025 : std_logic;
  signal gl_rom_n_1026, gl_rom_n_1027, gl_rom_n_1028, gl_rom_n_1029, gl_rom_n_1030 : std_logic;
  signal gl_rom_n_1031, gl_rom_n_1032, gl_rom_n_1033, gl_rom_n_1034, gl_rom_n_1035 : std_logic;
  signal gl_rom_n_1036, gl_rom_n_1037, gl_rom_n_1038, gl_rom_n_1039, gl_rom_n_1040 : std_logic;
  signal gl_rom_n_1041, gl_rom_n_1042, gl_rom_n_1043, gl_rom_n_1044, gl_rom_n_1045 : std_logic;
  signal gl_rom_n_1046, gl_rom_n_1047, gl_rom_n_1048, gl_rom_n_1049, gl_rom_n_1050 : std_logic;
  signal gl_rom_n_1051, gl_rom_n_1052, gl_rom_n_1053, gl_rom_n_1054, gl_rom_n_1055 : std_logic;
  signal gl_rom_n_1056, gl_rom_n_1057, gl_rom_n_1058, gl_rom_n_1059, gl_rom_n_1060 : std_logic;
  signal gl_rom_n_1061, gl_rom_n_1062, gl_rom_n_1063, gl_rom_n_1064, gl_rom_n_1065 : std_logic;
  signal gl_rom_n_1066, gl_rom_n_1067, gl_rom_n_1068, gl_rom_n_1069, gl_rom_n_1070 : std_logic;
  signal gl_rom_n_1071, gl_rom_n_1072, gl_rom_n_1073, gl_rom_n_1074, gl_rom_n_1075 : std_logic;
  signal gl_rom_n_1076, gl_rom_n_1077, gl_rom_n_1078, gl_rom_n_1079, gl_rom_n_1080 : std_logic;
  signal gl_rom_n_1081, gl_rom_n_1082, gl_rom_n_1083, gl_rom_n_1084, gl_rom_n_1085 : std_logic;
  signal gl_rom_n_1086, gl_rom_n_1087, gl_rom_n_1088, gl_rom_n_1089, gl_rom_n_1090 : std_logic;
  signal gl_rom_n_1091, gl_rom_n_1092, gl_rom_n_1093, gl_rom_n_1094, gl_rom_n_1095 : std_logic;
  signal gl_rom_n_1096, gl_rom_n_1097, gl_rom_n_1098, gl_rom_n_1099, gl_rom_n_1100 : std_logic;
  signal gl_rom_n_1101, gl_rom_n_1102, gl_rom_n_1103, gl_rom_n_1104, gl_rom_n_1105 : std_logic;
  signal gl_rom_n_1106, gl_rom_n_1107, gl_rom_n_1108, gl_rom_n_1109, gl_rom_n_1110 : std_logic;
  signal gl_rom_n_1111, gl_rom_n_1112, gl_rom_n_1113, gl_rom_n_1114, gl_rom_n_1115 : std_logic;
  signal gl_rom_n_1116, gl_rom_n_1117, gl_rom_n_1118, gl_rom_n_1119, gl_rom_n_1120 : std_logic;
  signal gl_rom_n_1121, gl_rom_n_1122, gl_rom_n_1123, gl_rom_n_1124, gl_rom_n_1125 : std_logic;
  signal gl_rom_n_1126, gl_rom_n_1127, gl_rom_n_1128, gl_rom_n_1129, gl_rom_n_1130 : std_logic;
  signal gl_rom_n_1131, gl_rom_n_1132, gl_rom_n_1133, gl_rom_n_1134, gl_rom_n_1135 : std_logic;
  signal gl_rom_n_1136, gl_rom_n_1137, gl_rom_n_1138, gl_rom_n_1139, gl_rom_n_1140 : std_logic;
  signal gl_rom_n_1141, gl_rom_n_1142, gl_rom_n_1143, gl_rom_n_1144, gl_rom_n_1145 : std_logic;
  signal gl_rom_n_1146, gl_rom_n_1147, gl_rom_n_1148, gl_rom_n_1149, gl_rom_n_1150 : std_logic;
  signal gl_rom_n_1151, gl_rom_n_1152, gl_rom_n_1153, gl_rom_n_1154, gl_rom_n_1155 : std_logic;
  signal gl_rom_n_1156, gl_rom_n_1157, gl_rom_n_1158, gl_rom_n_1159, gl_rom_n_1160 : std_logic;
  signal gl_rom_n_1161, gl_rom_n_1162, gl_rom_n_1163, gl_rom_n_1164, gl_rom_n_1165 : std_logic;
  signal gl_rom_n_1166, gl_rom_n_1167, gl_rom_n_1168, gl_rom_n_1169, gl_rom_n_1170 : std_logic;
  signal gl_rom_n_1171, gl_rom_n_1172, gl_rom_n_1173, gl_rom_n_1174, gl_rom_n_1175 : std_logic;
  signal gl_rom_n_1176, gl_rom_n_1177, gl_rom_n_1178, gl_rom_n_1179, gl_rom_n_1180 : std_logic;
  signal gl_rom_n_1181, gl_rom_n_1182, gl_rom_n_1183, gl_rom_n_1184, gl_rom_n_1185 : std_logic;
  signal gl_rom_n_1186, gl_rom_n_1187, gl_rom_n_1188, gl_rom_n_1189, gl_rom_n_1190 : std_logic;
  signal gl_rom_n_1191, gl_rom_n_1192, gl_rom_n_1193, gl_rom_n_1194, gl_rom_n_1195 : std_logic;
  signal gl_rom_n_1196, gl_rom_n_1197, gl_rom_n_1198, gl_rom_n_1199, gl_rom_n_1200 : std_logic;
  signal gl_rom_n_1201, gl_rom_n_1202, gl_rom_n_1203, gl_rom_n_1204, gl_rom_n_1205 : std_logic;
  signal gl_rom_n_1206, gl_rom_n_1207, gl_rom_n_1208, gl_rom_n_1209, gl_rom_n_1210 : std_logic;
  signal gl_rom_n_1211, gl_rom_n_1212, gl_rom_n_1213, gl_rom_n_1214, gl_rom_n_1215 : std_logic;
  signal gl_rom_n_1216, gl_rom_n_1217, gl_rom_n_1218, gl_rom_n_1219, gl_rom_n_1220 : std_logic;
  signal gl_rom_n_1221, gl_rom_n_1222, gl_rom_n_1223, gl_rom_n_1224, gl_rom_n_1225 : std_logic;
  signal gl_rom_n_1226, gl_rom_n_1227, gl_rom_n_1228, gl_rom_n_1229, gl_rom_n_1230 : std_logic;
  signal gl_rom_n_1231, gl_rom_n_1232, gl_rom_n_1233, gl_rom_n_1234, gl_rom_n_1235 : std_logic;
  signal gl_rom_n_1236, gl_rom_n_1237, gl_rom_n_1238, gl_rom_n_1239, gl_rom_n_1240 : std_logic;
  signal gl_rom_n_1241, gl_rom_n_1242, gl_rom_n_1243, gl_rom_n_1244, gl_rom_n_1245 : std_logic;
  signal gl_rom_n_1246, gl_rom_n_1247, gl_rom_n_1248, gl_rom_n_1249, gl_rom_n_1250 : std_logic;
  signal gl_rom_n_1251, gl_rom_n_1252, gl_rom_n_1253, gl_rom_n_1254, gl_rom_n_1255 : std_logic;
  signal gl_rom_n_1256, gl_rom_n_1257, gl_rom_n_1258, gl_rom_n_1259, gl_rom_n_1260 : std_logic;
  signal gl_rom_n_1261, gl_rom_n_1262, gl_rom_n_1263, gl_rom_n_1264, gl_rom_n_1265 : std_logic;
  signal gl_rom_n_1266, gl_rom_n_1267, gl_rom_n_1268, gl_rom_n_1269, gl_rom_n_1270 : std_logic;
  signal gl_rom_n_1271, gl_rom_n_1272, gl_rom_n_1273, gl_rom_n_1274, gl_rom_n_1275 : std_logic;
  signal gl_rom_n_1276, gl_rom_n_1277, gl_rom_n_1278, gl_rom_n_1279, gl_rom_n_1280 : std_logic;
  signal gl_rom_n_1281, gl_rom_n_1282, gl_rom_n_1283, gl_rom_n_1284, gl_rom_n_1285 : std_logic;
  signal gl_rom_n_1286, gl_rom_n_1287, gl_rom_n_1288, gl_rom_n_1289, gl_rom_n_1290 : std_logic;
  signal gl_rom_n_1291, gl_rom_n_1292, gl_rom_n_1293, gl_rom_n_1294, gl_rom_n_1295 : std_logic;
  signal gl_rom_n_1296, gl_rom_n_1297, gl_rom_n_1298, gl_rom_n_1299, gl_rom_n_1300 : std_logic;
  signal gl_rom_n_1301, gl_rom_n_1302, gl_rom_n_1303, gl_rom_n_1304, gl_rom_n_1305 : std_logic;
  signal gl_rom_n_1306, gl_rom_n_1307, gl_rom_n_1308, gl_rom_n_1309, gl_rom_n_1310 : std_logic;
  signal gl_rom_n_1311, gl_rom_n_1312, gl_rom_n_1313, gl_rom_n_1314, gl_rom_n_1315 : std_logic;
  signal gl_rom_n_1316, gl_rom_n_1317, gl_rom_n_1318, gl_rom_n_1319, gl_rom_n_1320 : std_logic;
  signal gl_rom_n_1321, gl_rom_n_1322, gl_rom_n_1323, gl_rom_n_1324, gl_rom_n_1325 : std_logic;
  signal gl_rom_n_1326, gl_rom_n_1327, gl_rom_n_1328, gl_rom_n_1329, gl_rom_n_1330 : std_logic;
  signal gl_rom_n_1331, gl_rom_n_1332, gl_rom_n_1333, gl_rom_n_1334, gl_rom_n_1335 : std_logic;
  signal gl_rom_n_1336, gl_rom_n_1337, gl_rom_n_1338, gl_rom_n_1339, gl_rom_n_1340 : std_logic;
  signal gl_rom_n_1341, gl_rom_n_1342, gl_rom_n_1343, gl_rom_n_1344, gl_rom_n_1345 : std_logic;
  signal gl_rom_n_1346, gl_rom_n_1347, gl_rom_n_1348, gl_rom_n_1349, gl_rom_n_1350 : std_logic;
  signal gl_rom_n_1351, gl_rom_n_1352, gl_rom_n_1353, gl_rom_n_1354, gl_rom_n_1355 : std_logic;
  signal gl_rom_n_1356, gl_rom_n_1357, gl_rom_n_1358, gl_rom_n_1359, gl_rom_n_1360 : std_logic;
  signal gl_rom_n_1361, gl_rom_n_1362, gl_rom_n_1363, gl_rom_n_1364, gl_rom_n_1365 : std_logic;
  signal gl_rom_n_1366, gl_rom_n_1367, gl_rom_n_1368, gl_rom_n_1369, gl_rom_n_1370 : std_logic;
  signal gl_rom_n_1371, gl_rom_n_1372, gl_rom_n_1373, gl_rom_n_1374, gl_rom_n_1375 : std_logic;
  signal gl_rom_n_1376, gl_rom_n_1377, gl_rom_n_1378, gl_rom_n_1379, gl_rom_n_1380 : std_logic;
  signal gl_rom_n_1381, gl_rom_n_1382, gl_rom_n_1383, gl_rom_n_1384, gl_rom_n_1385 : std_logic;
  signal gl_rom_n_1386, gl_rom_n_1387, gl_rom_n_1388, gl_rom_n_1389, gl_rom_n_1390 : std_logic;
  signal gl_rom_n_1391, gl_rom_n_1392, gl_rom_n_1393, gl_rom_n_1394, gl_rom_n_1395 : std_logic;
  signal gl_rom_n_1396, gl_rom_n_1397, gl_rom_n_1398, gl_rom_n_1399, gl_rom_n_1400 : std_logic;
  signal gl_rom_n_1401, gl_rom_n_1402, gl_rom_n_1403, gl_rom_n_1404, gl_rom_n_1405 : std_logic;
  signal gl_rom_n_1406, gl_rom_n_1407, gl_rom_n_1408, gl_rom_n_1409, gl_rom_n_1410 : std_logic;
  signal gl_rom_n_1411, gl_rom_n_1412, gl_rom_n_1413, gl_rom_n_1414, gl_rom_n_1415 : std_logic;
  signal gl_rom_n_1416, gl_rom_n_1417, gl_rom_n_1418, gl_rom_n_1419, gl_rom_n_1420 : std_logic;
  signal gl_rom_n_1421, gl_rom_n_1422, gl_rom_n_1423, gl_rom_n_1424, gl_rom_n_1425 : std_logic;
  signal gl_rom_n_1426, gl_rom_n_1427, gl_rom_n_1428, gl_rom_n_1429, gl_rom_n_1430 : std_logic;
  signal gl_rom_n_1431, gl_rom_n_1432, gl_rom_n_1433, gl_rom_n_1434, gl_rom_n_1435 : std_logic;
  signal gl_rom_n_1436, gl_rom_n_1437, gl_rom_n_1438, gl_rom_n_1439, gl_rom_n_1440 : std_logic;
  signal gl_rom_n_1441, gl_rom_n_1442, gl_rom_n_1443, gl_rom_n_1444, gl_rom_n_1445 : std_logic;
  signal gl_rom_n_1446, gl_rom_n_1447, gl_rom_n_1448, gl_rom_n_1449, gl_rom_n_1450 : std_logic;
  signal gl_rom_n_1451, gl_rom_n_1452, gl_rom_n_1453, gl_rom_n_1454, gl_rom_n_1455 : std_logic;
  signal gl_rom_n_1456, gl_rom_n_1457, gl_rom_n_1458, gl_rom_n_1459, gl_rom_n_1460 : std_logic;
  signal gl_rom_n_1461, gl_rom_n_1462, gl_rom_n_1463, gl_rom_n_1464, gl_rom_n_1465 : std_logic;
  signal gl_rom_n_1466, gl_rom_n_1467, gl_rom_n_1468, gl_rom_n_1469, gl_rom_n_1470 : std_logic;
  signal gl_rom_n_1471, gl_rom_n_1472, gl_rom_n_1473, gl_rom_n_1474, gl_rom_n_1475 : std_logic;
  signal gl_rom_n_1476, gl_rom_n_1477, gl_rom_n_1478, gl_rom_n_1479, gl_rom_n_1480 : std_logic;
  signal gl_rom_n_1481, gl_rom_n_1482, gl_rom_n_1483, gl_rom_n_1484, gl_rom_n_1485 : std_logic;
  signal gl_rom_n_1486, gl_rom_n_1487, gl_rom_n_1488, gl_rom_n_1489, gl_rom_n_1490 : std_logic;
  signal gl_rom_n_1491, gl_rom_n_1492, gl_rom_n_1493, gl_rom_n_1494, gl_rom_n_1495 : std_logic;
  signal gl_rom_n_1496, gl_rom_n_1497, gl_rom_n_1498, gl_rom_n_1499, gl_rom_n_1500 : std_logic;
  signal gl_sig_blue, gl_sig_green, gl_sig_red, gl_sig_scale_h, gl_sig_scale_v : std_logic;
  signal gl_sig_v, gl_vga_buf_Bint, gl_vga_buf_Gint, gl_vga_buf_Hint, gl_vga_buf_Rint : std_logic;
  signal gl_vga_buf_Vint, gl_vgd_n_0, gl_vgd_n_2, gl_vgd_n_3, gl_vgd_n_4 : std_logic;
  signal gl_vgd_n_5, gl_vgd_n_6, gl_vgd_n_7, gl_vgd_n_8, gl_vgd_n_9 : std_logic;
  signal gl_vgd_n_10, gl_vgd_n_11, gl_vgd_n_12, gl_vgd_n_13, gl_vgd_n_14 : std_logic;
  signal gl_vgd_n_15, gl_vgd_n_16, gl_vgd_n_17, gl_vgd_n_18, gl_vgd_n_19 : std_logic;
  signal gl_vgd_n_20, gl_vgd_n_21, gl_vgd_n_22, gl_vgd_n_23, gl_vgd_n_24 : std_logic;
  signal gl_vgd_n_25, gl_vgd_n_26, gl_vgd_n_27, gl_vgd_n_28, gl_vgd_n_29 : std_logic;
  signal gl_vgd_n_30, gl_vgd_n_31, gl_vgd_n_32, gl_vgd_n_33, gl_vgd_n_34 : std_logic;
  signal gl_vgd_n_35, gl_vgd_n_36, gl_vgd_n_37, gl_vgd_n_38, gl_vgd_n_39 : std_logic;
  signal gl_vgd_n_40, gl_vgd_n_41, gl_vgd_n_42, gl_vgd_n_43, gl_vgd_n_44 : std_logic;
  signal gl_vgd_n_45, gl_vgd_n_46, gl_vgd_n_47, gl_vgd_n_48, gl_vgd_n_49 : std_logic;
  signal gl_vgd_n_50, gl_vgd_n_51, gl_vgd_n_52, gl_vgd_n_53, gl_vgd_n_54 : std_logic;
  signal gl_vgd_n_55, gl_vgd_n_56, gl_vgd_n_57, gl_vgd_n_58, gl_vgd_n_59 : std_logic;
  signal gl_vgd_n_60, gl_vgd_n_61, gl_vgd_n_62, gl_vgd_n_63, gl_vgd_n_64 : std_logic;
  signal gl_vgd_n_65, gl_vgd_n_67, gl_vgd_n_68, gl_vgd_n_69, gl_vgd_n_70 : std_logic;
  signal gl_vgd_n_71, gl_vgd_n_72, gl_vgd_n_73, gl_vgd_n_74, gl_vgd_n_75 : std_logic;
  signal gl_vgd_n_76, gl_vgd_n_77, gl_vgd_n_78, gl_vgd_n_79, gl_vgd_n_80 : std_logic;
  signal ml_handshake_mouse_out, ml_il_color1_n_0, ml_il_color1_n_1, ml_il_color1_n_3, ml_il_color1_n_4 : std_logic;
  signal ml_il_color1_n_5, ml_il_color1_n_6, ml_il_color1_n_7, ml_il_color1_n_8, ml_il_color1_n_9 : std_logic;
  signal ml_il_color1_n_10, ml_il_color1_n_11, ml_il_color1_n_12, ml_il_color1_n_13, ml_il_color1_n_14 : std_logic;
  signal ml_il_color1_n_15, ml_il_color1_n_16, ml_il_color1_n_17, ml_il_color1_n_18, ml_il_color1_n_23 : std_logic;
  signal ml_il_color1_n_24, ml_il_x1_n_1, ml_il_x1_n_2, ml_il_x1_n_5, ml_il_x1_n_6 : std_logic;
  signal ml_il_x1_n_7, ml_il_x1_n_8, ml_il_x1_n_9, ml_il_x1_n_10, ml_il_x1_n_11 : std_logic;
  signal ml_il_x1_n_12, ml_il_x1_n_13, ml_il_x1_n_14, ml_il_x1_n_15, ml_il_x1_n_16 : std_logic;
  signal ml_il_x1_n_17, ml_il_x1_n_18, ml_il_x1_n_19, ml_il_x1_n_20, ml_il_x1_n_21 : std_logic;
  signal ml_il_x1_n_22, ml_il_x1_n_23, ml_il_x1_n_24, ml_il_x1_n_25, ml_il_x1_n_26 : std_logic;
  signal ml_il_x1_n_27, ml_il_x1_n_28, ml_il_x1_n_43, ml_il_x1_n_44, ml_il_x1_n_46 : std_logic;
  signal ml_il_x1_n_47, ml_il_x1_n_48, ml_il_x1_n_49, ml_il_x1_n_50, ml_il_x1_n_51 : std_logic;
  signal ml_il_x1_n_52, ml_il_y1_n_1, ml_il_y1_n_2, ml_il_y1_n_5, ml_il_y1_n_6 : std_logic;
  signal ml_il_y1_n_7, ml_il_y1_n_8, ml_il_y1_n_9, ml_il_y1_n_10, ml_il_y1_n_11 : std_logic;
  signal ml_il_y1_n_12, ml_il_y1_n_13, ml_il_y1_n_14, ml_il_y1_n_15, ml_il_y1_n_16 : std_logic;
  signal ml_il_y1_n_17, ml_il_y1_n_18, ml_il_y1_n_19, ml_il_y1_n_20, ml_il_y1_n_21 : std_logic;
  signal ml_il_y1_n_22, ml_il_y1_n_23, ml_il_y1_n_24, ml_il_y1_n_25, ml_il_y1_n_26 : std_logic;
  signal ml_il_y1_n_27, ml_il_y1_n_28, ml_il_y1_n_43, ml_il_y1_n_44, ml_il_y1_n_46 : std_logic;
  signal ml_il_y1_n_47, ml_il_y1_n_48, ml_il_y1_n_49, ml_il_y1_n_50, ml_il_y1_n_51 : std_logic;
  signal ml_il_y1_n_52, ml_ms_actBit, ml_ms_btnflipfloprst, ml_ms_cntD_n_0, ml_ms_cntD_n_1 : std_logic;
  signal ml_ms_cntD_n_2, ml_ms_cntD_n_3, ml_ms_cntD_n_4, ml_ms_cntD_n_5, ml_ms_cntD_n_6 : std_logic;
  signal ml_ms_cntD_n_7, ml_ms_cntD_n_8, ml_ms_cntD_n_9, ml_ms_cntD_n_10, ml_ms_cntD_n_11 : std_logic;
  signal ml_ms_cntD_n_12, ml_ms_cntD_n_13, ml_ms_cntD_n_14, ml_ms_cntD_n_15, ml_ms_cntD_n_16 : std_logic;
  signal ml_ms_cntD_n_17, ml_ms_cntD_n_18, ml_ms_cntD_n_19, ml_ms_cntD_n_20, ml_ms_cntD_n_21 : std_logic;
  signal ml_ms_cntD_n_22, ml_ms_cntD_n_23, ml_ms_cntReset15K, ml_ms_cntReset25M, ml_ms_cntReset25M_main : std_logic;
  signal ml_ms_cntReset25M_send, ml_ms_cnt_n_0, ml_ms_cnt_n_1, ml_ms_cnt_n_2, ml_ms_cnt_n_3 : std_logic;
  signal ml_ms_cnt_n_4, ml_ms_cnt_n_5, ml_ms_cnt_n_6, ml_ms_cnt_n_7, ml_ms_cnt_n_8 : std_logic;
  signal ml_ms_cnt_n_9, ml_ms_cnt_n_10, ml_ms_cnt_n_11, ml_ms_cnt_n_12, ml_ms_cnt_n_13 : std_logic;
  signal ml_ms_cnt_n_14, ml_ms_cnt_n_15, ml_ms_cnt_n_16, ml_ms_cnt_n_17, ml_ms_cnt_n_18 : std_logic;
  signal ml_ms_cnt_n_19, ml_ms_cnt_n_20, ml_ms_cnt_n_21, ml_ms_cnt_n_22, ml_ms_cnt_n_23 : std_logic;
  signal ml_ms_count_debounce_reset, ml_ms_ed_n_0, ml_ms_ed_n_1, ml_ms_ed_n_2, ml_ms_ed_n_3 : std_logic;
  signal ml_ms_ed_n_4, ml_ms_ed_n_5, ml_ms_ed_n_6, ml_ms_ed_n_7, ml_ms_ed_n_8 : std_logic;
  signal ml_ms_ed_n_9, ml_ms_ed_reg1, ml_ms_ed_reg2, ml_ms_mfsm_n_0, ml_ms_mfsm_n_1 : std_logic;
  signal ml_ms_mfsm_n_3, ml_ms_mfsm_n_4, ml_ms_mfsm_n_5, ml_ms_mfsm_n_6, ml_ms_mfsm_n_7 : std_logic;
  signal ml_ms_mfsm_n_8, ml_ms_mfsm_n_9, ml_ms_mfsm_n_10, ml_ms_mfsm_n_11, ml_ms_mfsm_n_12 : std_logic;
  signal ml_ms_mfsm_n_13, ml_ms_mfsm_n_14, ml_ms_mfsm_n_15, ml_ms_mfsm_n_16, ml_ms_mfsm_n_17 : std_logic;
  signal ml_ms_mfsm_n_18, ml_ms_mfsm_n_19, ml_ms_mfsm_n_20, ml_ms_mfsm_n_21, ml_ms_mfsm_n_22 : std_logic;
  signal ml_ms_mfsm_n_23, ml_ms_mfsm_n_24, ml_ms_mfsm_n_25, ml_ms_mfsm_n_26, ml_ms_mfsm_n_27 : std_logic;
  signal ml_ms_mfsm_n_28, ml_ms_mfsm_n_29, ml_ms_mfsm_n_30, ml_ms_mfsm_n_31, ml_ms_mfsm_n_32 : std_logic;
  signal ml_ms_mfsm_n_33, ml_ms_mfsm_n_34, ml_ms_mfsm_n_35, ml_ms_mfsm_n_36, ml_ms_mfsm_n_37 : std_logic;
  signal ml_ms_mfsm_n_38, ml_ms_mfsm_n_39, ml_ms_mfsm_n_40, ml_ms_mfsm_n_41, ml_ms_mfsm_n_42 : std_logic;
  signal ml_ms_mfsm_n_43, ml_ms_mfsm_n_44, ml_ms_mfsm_n_45, ml_ms_mfsm_n_46, ml_ms_mfsm_n_47 : std_logic;
  signal ml_ms_mfsm_n_48, ml_ms_mfsm_n_49, ml_ms_mfsm_n_50, ml_ms_mfsm_n_51, ml_ms_mfsm_n_52 : std_logic;
  signal ml_ms_mfsm_n_53, ml_ms_mfsm_n_54, ml_ms_mfsm_n_55, ml_ms_mfsm_n_56, ml_ms_mfsm_n_57 : std_logic;
  signal ml_ms_mfsm_n_58, ml_ms_mfsm_n_59, ml_ms_mfsm_n_60, ml_ms_mfsm_n_61, ml_ms_mfsm_n_62 : std_logic;
  signal ml_ms_mfsm_n_63, ml_ms_mfsm_n_64, ml_ms_mfsm_n_66, ml_ms_mfsm_n_116, ml_ms_mfsm_n_117 : std_logic;
  signal ml_ms_mfsm_n_118, ml_ms_muxFSM, ml_ms_muxReg, ml_ms_mux_select, ml_ms_mux_select_main : std_logic;
  signal ml_ms_mx_n_0, ml_ms_mx_n_1, ml_ms_n_0, ml_ms_n_1, ml_ms_n_2 : std_logic;
  signal ml_ms_n_3, ml_ms_n_4, ml_ms_n_5, ml_ms_n_6, ml_ms_n_7 : std_logic;
  signal ml_ms_n_8, ml_ms_n_9, ml_ms_n_10, ml_ms_n_11, ml_ms_n_12 : std_logic;
  signal ml_ms_n_13, ml_ms_n_14, ml_ms_n_15, ml_ms_n_16, ml_ms_n_17 : std_logic;
  signal ml_ms_n_18, ml_ms_n_19, ml_ms_n_20, ml_ms_n_21, ml_ms_n_22 : std_logic;
  signal ml_ms_n_23, ml_ms_n_24, ml_ms_n_25, ml_ms_n_26, ml_ms_n_27 : std_logic;
  signal ml_ms_n_28, ml_ms_n_29, ml_ms_n_30, ml_ms_n_31, ml_ms_n_32 : std_logic;
  signal ml_ms_n_33, ml_ms_n_34, ml_ms_n_35, ml_ms_n_36, ml_ms_n_37 : std_logic;
  signal ml_ms_n_38, ml_ms_n_39, ml_ms_n_40, ml_ms_n_41, ml_ms_n_42 : std_logic;
  signal ml_ms_n_43, ml_ms_n_44, ml_ms_n_45, ml_ms_n_46, ml_ms_n_47 : std_logic;
  signal ml_ms_n_48, ml_ms_n_49, ml_ms_n_50, ml_ms_n_51, ml_ms_n_52 : std_logic;
  signal ml_ms_n_53, ml_ms_n_54, ml_ms_n_55, ml_ms_n_56, ml_ms_n_57 : std_logic;
  signal ml_ms_n_58, ml_ms_n_59, ml_ms_n_60, ml_ms_n_61, ml_ms_n_62 : std_logic;
  signal ml_ms_n_63, ml_ms_output_edgedet, ml_ms_reset_send, ml_ms_sfsm_n_383, ml_ms_sr11_data_out_0_79 : std_logic;
  signal ml_ms_sr11_data_out_1_80, ml_ms_sr11_data_out_5_84, ml_ms_tb_n_0, ml_ms_tb_n_1, ml_ms_tb_n_2 : std_logic;
  signal ml_ms_tb_n_3, ml_ms_tb_n_4, ml_ms_tb_n_5, ml_ms_tb_n_6, ml_ms_xflipfloprst : std_logic;
  signal ml_ms_yflipfloprst, sig_countlow, sig_draw, sig_middelsteknop, sig_rescount : std_logic;

begin

  FE_PHC672_gl_ram_n_470 : BUFFD1P5BWP7T port map(I => gl_ram_n_470, Z => FE_PHN672_gl_ram_n_470);
  FE_PHC671_gl_ram_n_435 : DEL01BWP7T port map(I => gl_ram_n_435, Z => FE_PHN671_gl_ram_n_435);
  FE_PHC670_gl_ram_ram_35_0 : DEL01BWP7T port map(I => FE_PHN583_gl_ram_ram_35_0, Z => FE_PHN670_gl_ram_ram_35_0);
  FE_PHC669_gl_ram_ram_27_2 : BUFFD1P5BWP7T port map(I => FE_PHN669_gl_ram_ram_27_2, Z => gl_ram_ram_27(2));
  FE_PHC668_gl_ram_ram_1_2 : DEL02BWP7T port map(I => FE_PHN519_gl_ram_ram_1_2, Z => FE_PHN668_gl_ram_ram_1_2);
  FE_PHC667_gl_ram_ram_33_0 : DEL01BWP7T port map(I => gl_ram_ram_33(0), Z => FE_PHN667_gl_ram_ram_33_0);
  FE_PHC666_ml_ms_count_debounce_12 : DEL01BWP7T port map(I => FE_PHN653_ml_ms_count_debounce_12, Z => FE_PHN666_ml_ms_count_debounce_12);
  FE_PHC665_gl_ram_ram_21_0 : DEL01BWP7T port map(I => FE_PHN522_gl_ram_ram_21_0, Z => FE_PHN665_gl_ram_ram_21_0);
  FE_PHC664_gl_ram_ram_58_1 : DEL01BWP7T port map(I => FE_PHN664_gl_ram_ram_58_1, Z => gl_ram_ram_58(1));
  FE_PHC663_ml_ms_count_debounce_12 : BUFFD3BWP7T port map(I => FE_PHN615_ml_ms_count_debounce_12, Z => FE_PHN663_ml_ms_count_debounce_12);
  FE_PHC662_gl_ram_ram_37_2 : BUFFD3BWP7T port map(I => FE_PHN593_gl_ram_ram_37_2, Z => FE_PHN662_gl_ram_ram_37_2);
  FE_PHC661_gl_ram_ram_75_0 : DEL01BWP7T port map(I => FE_PHN661_gl_ram_ram_75_0, Z => gl_ram_ram_75(0));
  FE_PHC660_gl_ram_ram_59_2 : DEL02BWP7T port map(I => FE_PHN660_gl_ram_ram_59_2, Z => gl_ram_ram_59(2));
  FE_PHC659_gl_ram_ram_18_0 : BUFFD1P5BWP7T port map(I => FE_PHN599_gl_ram_ram_18_0, Z => FE_PHN659_gl_ram_ram_18_0);
  FE_PHC658_gl_ram_ram_43_1 : CKBD0BWP7T port map(I => gl_ram_ram_43(1), Z => FE_PHN658_gl_ram_ram_43_1);
  FE_PHC657_gl_ram_n_445 : CKBD0BWP7T port map(I => gl_ram_n_445, Z => FE_PHN657_gl_ram_n_445);
  FE_PHC656_ml_ms_ed_n_8 : CKBD0BWP7T port map(I => FE_PHN551_ml_ms_ed_n_8, Z => FE_PHN656_ml_ms_ed_n_8);
  FE_PHC655_ml_ms_count_debounce_7 : DEL01BWP7T port map(I => FE_PHN612_ml_ms_count_debounce_7, Z => FE_PHN655_ml_ms_count_debounce_7);
  FE_PHC654_gl_ram_ram_17_1 : DEL01BWP7T port map(I => gl_ram_ram_17(1), Z => FE_PHN654_gl_ram_ram_17_1);
  FE_PHC653_ml_ms_count_debounce_12 : CKBD0BWP7T port map(I => FE_PHN615_ml_ms_count_debounce_12, Z => FE_PHN653_ml_ms_count_debounce_12);
  FE_PHC652_gl_ram_ram_11_2 : BUFFD1P5BWP7T port map(I => FE_PHN652_gl_ram_ram_11_2, Z => gl_ram_ram_11(2));
  FE_PHC651_gl_ram_ram_16_2 : DEL01BWP7T port map(I => FE_PHN651_gl_ram_ram_16_2, Z => gl_ram_ram_16(2));
  FE_PHC650_gl_ram_ram_97_1 : BUFFD3BWP7T port map(I => FE_PHN608_gl_ram_ram_97_1, Z => FE_PHN650_gl_ram_ram_97_1);
  FE_PHC649_gl_ram_ram_34_1 : DEL01BWP7T port map(I => gl_ram_ram_34(1), Z => FE_PHN649_gl_ram_ram_34_1);
  FE_PHC648_gl_ram_ram_9_2 : BUFFD1P5BWP7T port map(I => FE_PHN528_gl_ram_ram_9_2, Z => FE_PHN648_gl_ram_ram_9_2);
  FE_PHC647_gl_ram_ram_8_1 : DEL01BWP7T port map(I => FE_PHN647_gl_ram_ram_8_1, Z => gl_ram_ram_8(1));
  FE_PHC646_gl_ram_ram_8_2 : BUFFD1P5BWP7T port map(I => gl_ram_ram_8(2), Z => FE_PHN646_gl_ram_ram_8_2);
  FE_PHC645_gl_ram_ram_51_2 : BUFFD2BWP7T port map(I => gl_ram_ram_51(2), Z => FE_PHN645_gl_ram_ram_51_2);
  FE_PHC644_gl_ram_ram_12_2 : DEL01BWP7T port map(I => FE_PHN607_gl_ram_ram_12_2, Z => FE_PHN644_gl_ram_ram_12_2);
  FE_PHC643_gl_ram_ram_88_0 : DEL01BWP7T port map(I => gl_ram_ram_88(0), Z => FE_PHN643_gl_ram_ram_88_0);
  FE_PHC642_gl_ram_ram_12_1 : CKBD0BWP7T port map(I => FE_PHN642_gl_ram_ram_12_1, Z => gl_ram_ram_12(1));
  FE_PHC641_ml_ms_sr_new_new_data_4 : DEL01BWP7T port map(I => ml_ms_sr_new_new_data(4), Z => FE_PHN641_ml_ms_sr_new_new_data_4);
  FE_PHC640_gl_ram_ram_91_1 : BUFFD1P5BWP7T port map(I => gl_ram_ram_91(1), Z => FE_PHN640_gl_ram_ram_91_1);
  FE_PHC639_gl_ram_ram_27_0 : DEL01BWP7T port map(I => gl_ram_ram_27(0), Z => FE_PHN639_gl_ram_ram_27_0);
  FE_PHC638_gl_ram_ram_5_1 : DEL01BWP7T port map(I => gl_ram_ram_5(1), Z => FE_PHN638_gl_ram_ram_5_1);
  FE_PHC637_gl_ram_ram_48_1 : DEL01BWP7T port map(I => FE_PHN584_gl_ram_ram_48_1, Z => FE_PHN637_gl_ram_ram_48_1);
  FE_PHC636_ml_ms_ed_reg2 : DEL01BWP7T port map(I => ml_ms_ed_reg2, Z => FE_PHN636_ml_ms_ed_reg2);
  FE_PHC635_gl_ram_ram_27_2 : DEL02BWP7T port map(I => FE_PHN518_gl_ram_ram_27_2, Z => FE_PHN635_gl_ram_ram_27_2);
  FE_PHC634_gl_ram_ram_50_2 : BUFFD1P5BWP7T port map(I => FE_PHN589_gl_ram_ram_50_2, Z => FE_PHN634_gl_ram_ram_50_2);
  FE_PHC633_gl_ram_ram_50_1 : BUFFD1P5BWP7T port map(I => FE_PHN588_gl_ram_ram_50_1, Z => FE_PHN633_gl_ram_ram_50_1);
  FE_PHC632_gl_ram_ram_57_1 : DEL01BWP7T port map(I => FE_PHN581_gl_ram_ram_57_1, Z => FE_PHN632_gl_ram_ram_57_1);
  FE_PHC631_gl_ram_ram_33_2 : DEL01BWP7T port map(I => gl_ram_ram_33(2), Z => FE_PHN631_gl_ram_ram_33_2);
  FE_PHC630_gl_ram_ram_25_0 : DEL01BWP7T port map(I => FE_PHN577_gl_ram_ram_25_0, Z => FE_PHN630_gl_ram_ram_25_0);
  FE_PHC629_gl_ram_ram_29_1 : DEL01BWP7T port map(I => FE_PHN587_gl_ram_ram_29_1, Z => FE_PHN629_gl_ram_ram_29_1);
  FE_PHC628_gl_ram_n_437 : CKBD0BWP7T port map(I => gl_ram_n_437, Z => FE_PHN628_gl_ram_n_437);
  FE_PHC627_gl_ram_n_523 : DEL01BWP7T port map(I => gl_ram_n_523, Z => FE_PHN627_gl_ram_n_523);
  FE_PHC626_gl_ram_ram_41_0 : CKBD0BWP7T port map(I => gl_ram_ram_41(0), Z => FE_PHN626_gl_ram_ram_41_0);
  FE_PHC625_gl_ram_ram_4_0 : DEL01BWP7T port map(I => FE_PHN603_gl_ram_ram_4_0, Z => FE_PHN625_gl_ram_ram_4_0);
  FE_PHC624_gl_ram_ram_89_0 : DEL01BWP7T port map(I => FE_PHN594_gl_ram_ram_89_0, Z => FE_PHN624_gl_ram_ram_89_0);
  FE_PHC623_ml_ms_sr_new_new_data_0 : DEL01BWP7T port map(I => FE_PHN613_ml_ms_sr_new_new_data_0, Z => FE_PHN623_ml_ms_sr_new_new_data_0);
  FE_PHC622_ml_ms_ed_n_8 : CKBD0BWP7T port map(I => FE_PHN656_ml_ms_ed_n_8, Z => FE_PHN622_ml_ms_ed_n_8);
  FE_PHC621_ml_ms_ed_n_2 : CKBD2BWP7T port map(I => FE_PHN470_ml_ms_ed_n_2, Z => FE_PHN621_ml_ms_ed_n_2);
  FE_PHC620_ml_ms_n_23 : DEL01BWP7T port map(I => FE_PHN620_ml_ms_n_23, Z => ml_ms_n_23);
  FE_PHC619_ml_ms_n_24 : CKBD0BWP7T port map(I => FE_PHN459_ml_ms_n_24, Z => FE_PHN619_ml_ms_n_24);
  FE_PHC618_ml_ms_n_22 : CKBD0BWP7T port map(I => ml_ms_n_22, Z => FE_PHN618_ml_ms_n_22);
  FE_PHC617_ml_ms_count_debounce_10 : DEL01BWP7T port map(I => FE_PHN463_ml_ms_count_debounce_10, Z => FE_PHN617_ml_ms_count_debounce_10);
  FE_PHC616_ml_ms_count_debounce_6 : DEL01BWP7T port map(I => ml_ms_count_debounce(6), Z => FE_PHN616_ml_ms_count_debounce_6);
  FE_PHC615_ml_ms_count_debounce_12 : BUFFD1P5BWP7T port map(I => ml_ms_count_debounce(12), Z => FE_PHN615_ml_ms_count_debounce_12);
  FE_PHC614_ml_ms_ed_state_0 : DEL02BWP7T port map(I => FE_PHN614_ml_ms_ed_state_0, Z => ml_ms_ed_state(0));
  FE_PHC613_ml_ms_sr_new_new_data_0 : CKBD0BWP7T port map(I => ml_ms_sr_new_new_data(0), Z => FE_PHN613_ml_ms_sr_new_new_data_0);
  FE_PHC612_ml_ms_count_debounce_7 : CKBD0BWP7T port map(I => ml_ms_count_debounce(7), Z => FE_PHN612_ml_ms_count_debounce_7);
  FE_PHC611_gl_ram_ram_19_1 : DEL015BWP7T port map(I => FE_PHN611_gl_ram_ram_19_1, Z => gl_ram_ram_19(1));
  FE_PHC610_ml_ms_ed_state_1 : DEL02BWP7T port map(I => ml_ms_ed_state(1), Z => FE_PHN610_ml_ms_ed_state_1);
  FE_PHC609_gl_ram_ram_17_1 : CKBD0BWP7T port map(I => FE_PHN654_gl_ram_ram_17_1, Z => FE_PHN609_gl_ram_ram_17_1);
  FE_PHC608_gl_ram_ram_97_1 : CKBD2BWP7T port map(I => FE_PHN480_gl_ram_ram_97_1, Z => FE_PHN608_gl_ram_ram_97_1);
  FE_PHC607_gl_ram_ram_12_2 : CKBD2BWP7T port map(I => FE_PHN535_gl_ram_ram_12_2, Z => FE_PHN607_gl_ram_ram_12_2);
  FE_PHC606_gl_ram_ram_58_1 : DEL02BWP7T port map(I => FE_PHN520_gl_ram_ram_58_1, Z => FE_PHN606_gl_ram_ram_58_1);
  FE_PHC605_gl_ram_ram_24_2 : DEL02BWP7T port map(I => FE_PHN521_gl_ram_ram_24_2, Z => FE_PHN605_gl_ram_ram_24_2);
  FE_PHC604_gl_ram_ram_73_2 : BUFFD1P5BWP7T port map(I => FE_PHN472_gl_ram_ram_73_2, Z => FE_PHN604_gl_ram_ram_73_2);
  FE_PHC603_gl_ram_ram_4_0 : BUFFD0BWP7T port map(I => gl_ram_ram_4(0), Z => FE_PHN603_gl_ram_ram_4_0);
  FE_PHC602_gl_ram_ram_88_0 : CKBD0BWP7T port map(I => FE_PHN514_gl_ram_ram_88_0, Z => FE_PHN602_gl_ram_ram_88_0);
  FE_PHC601_gl_ram_ram_21_0 : DEL02BWP7T port map(I => FE_PHN665_gl_ram_ram_21_0, Z => FE_PHN601_gl_ram_ram_21_0);
  FE_PHC600_gl_ram_ram_32_1 : CKBD0BWP7T port map(I => FE_PHN497_gl_ram_ram_32_1, Z => FE_PHN600_gl_ram_ram_32_1);
  FE_PHC599_gl_ram_ram_18_0 : CKBD0BWP7T port map(I => gl_ram_ram_18(0), Z => FE_PHN599_gl_ram_ram_18_0);
  FE_PHC598_gl_ram_ram_16_2 : CKBD0BWP7T port map(I => gl_ram_ram_16(2), Z => FE_PHN598_gl_ram_ram_16_2);
  FE_PHC597_gl_ram_ram_2_2 : DEL015BWP7T port map(I => FE_PHN517_gl_ram_ram_2_2, Z => FE_PHN597_gl_ram_ram_2_2);
  FE_PHC596_gl_ram_ram_27_0 : CKBD0BWP7T port map(I => FE_PHN530_gl_ram_ram_27_0, Z => FE_PHN596_gl_ram_ram_27_0);
  FE_PHC595_gl_ram_ram_12_1 : CKBD0BWP7T port map(I => FE_PHN504_gl_ram_ram_12_1, Z => FE_PHN595_gl_ram_ram_12_1);
  FE_PHC594_gl_ram_ram_89_0 : CKBD0BWP7T port map(I => FE_PHN531_gl_ram_ram_89_0, Z => FE_PHN594_gl_ram_ram_89_0);
  FE_PHC593_gl_ram_ram_37_2 : BUFFD1P5BWP7T port map(I => FE_PHN509_gl_ram_ram_37_2, Z => FE_PHN593_gl_ram_ram_37_2);
  FE_PHC592_gl_ram_ram_35_2 : CKBD0BWP7T port map(I => FE_PHN477_gl_ram_ram_35_2, Z => FE_PHN592_gl_ram_ram_35_2);
  FE_PHC591_gl_ram_ram_56_2 : CKBD0BWP7T port map(I => FE_PHN500_gl_ram_ram_56_2, Z => FE_PHN591_gl_ram_ram_56_2);
  FE_PHC590_gl_ram_ram_56_1 : CKBD0BWP7T port map(I => FE_PHN501_gl_ram_ram_56_1, Z => FE_PHN590_gl_ram_ram_56_1);
  FE_PHC589_gl_ram_ram_50_2 : CKBD0BWP7T port map(I => FE_PHN537_gl_ram_ram_50_2, Z => FE_PHN589_gl_ram_ram_50_2);
  FE_PHC588_gl_ram_ram_50_1 : CKBD0BWP7T port map(I => FE_PHN474_gl_ram_ram_50_1, Z => FE_PHN588_gl_ram_ram_50_1);
  FE_PHC587_gl_ram_ram_29_1 : CKBD0BWP7T port map(I => FE_PHN495_gl_ram_ram_29_1, Z => FE_PHN587_gl_ram_ram_29_1);
  FE_PHC586_gl_ram_ram_51_2 : CKBD0BWP7T port map(I => FE_PHN502_gl_ram_ram_51_2, Z => FE_PHN586_gl_ram_ram_51_2);
  FE_PHC585_gl_ram_ram_33_0 : CKBD0BWP7T port map(I => FE_PHN488_gl_ram_ram_33_0, Z => FE_PHN585_gl_ram_ram_33_0);
  FE_PHC584_gl_ram_ram_48_1 : CKBD0BWP7T port map(I => FE_PHN490_gl_ram_ram_48_1, Z => FE_PHN584_gl_ram_ram_48_1);
  FE_PHC583_gl_ram_ram_35_0 : CKBD0BWP7T port map(I => FE_PHN493_gl_ram_ram_35_0, Z => FE_PHN583_gl_ram_ram_35_0);
  FE_PHC582_gl_ram_ram_41_0 : CKBD0BWP7T port map(I => FE_PHN536_gl_ram_ram_41_0, Z => FE_PHN582_gl_ram_ram_41_0);
  FE_PHC581_gl_ram_ram_57_1 : CKBD0BWP7T port map(I => FE_PHN539_gl_ram_ram_57_1, Z => FE_PHN581_gl_ram_ram_57_1);
  FE_PHC580_gl_ram_ram_75_0 : CKBD0BWP7T port map(I => FE_PHN498_gl_ram_ram_75_0, Z => FE_PHN580_gl_ram_ram_75_0);
  FE_PHC579_gl_ram_n_489 : DEL02BWP7T port map(I => FE_PHN579_gl_ram_n_489, Z => gl_ram_n_489);
  FE_PHC578_gl_ram_ram_8_2 : CKBD0BWP7T port map(I => FE_PHN541_gl_ram_ram_8_2, Z => FE_PHN578_gl_ram_ram_8_2);
  FE_PHC577_gl_ram_ram_25_0 : CKBD0BWP7T port map(I => FE_PHN540_gl_ram_ram_25_0, Z => FE_PHN577_gl_ram_ram_25_0);
  FE_PHC576_gl_ram_ram_33_2 : CKBD0BWP7T port map(I => FE_PHN482_gl_ram_ram_33_2, Z => FE_PHN576_gl_ram_ram_33_2);
  FE_PHC575_gl_ram_ram_8_0 : CKBD0BWP7T port map(I => FE_PHN499_gl_ram_ram_8_0, Z => FE_PHN575_gl_ram_ram_8_0);
  FE_PHC574_gl_ram_ram_91_1 : CKBD0BWP7T port map(I => FE_PHN479_gl_ram_ram_91_1, Z => FE_PHN574_gl_ram_ram_91_1);
  FE_PHC573_gl_ram_ram_11_2 : CKBD0BWP7T port map(I => gl_ram_ram_11(2), Z => FE_PHN573_gl_ram_ram_11_2);
  FE_PHC572_gl_ram_ram_8_1 : CKBD0BWP7T port map(I => FE_PHN534_gl_ram_ram_8_1, Z => FE_PHN572_gl_ram_ram_8_1);
  FE_PHC571_gl_ram_ram_34_1 : CKBD0BWP7T port map(I => FE_PHN475_gl_ram_ram_34_1, Z => FE_PHN571_gl_ram_ram_34_1);
  FE_PHC570_gl_ram_ram_82_0 : DEL01BWP7T port map(I => FE_PHN462_gl_ram_ram_82_0, Z => FE_PHN570_gl_ram_ram_82_0);
  FE_PHC569_gl_ram_ram_2_0 : BUFFD3BWP7T port map(I => FE_PHN505_gl_ram_ram_2_0, Z => FE_PHN569_gl_ram_ram_2_0);
  FE_PHC568_gl_ram_ram_11_1 : BUFFD3BWP7T port map(I => FE_PHN508_gl_ram_ram_11_1, Z => FE_PHN568_gl_ram_ram_11_1);
  FE_PHC567_gl_ram_ram_3_2 : BUFFD3BWP7T port map(I => FE_PHN503_gl_ram_ram_3_2, Z => FE_PHN567_gl_ram_ram_3_2);
  FE_PHC566_ml_ms_muxReg : BUFFD0BWP7T port map(I => ml_ms_muxReg, Z => FE_PHN566_ml_ms_muxReg);
  FE_PHC565_gl_ram_ram_9_0 : BUFFD3BWP7T port map(I => FE_PHN491_gl_ram_ram_9_0, Z => FE_PHN565_gl_ram_ram_9_0);
  FE_PHC564_gl_ram_ram_43_2 : BUFFD2BWP7T port map(I => FE_PHN512_gl_ram_ram_43_2, Z => FE_PHN564_gl_ram_ram_43_2);
  FE_PHC563_gl_ram_ram_24_0 : BUFFD3BWP7T port map(I => FE_PHN496_gl_ram_ram_24_0, Z => FE_PHN563_gl_ram_ram_24_0);
  FE_PHC562_gl_ram_ram_3_0 : BUFFD3BWP7T port map(I => FE_PHN487_gl_ram_ram_3_0, Z => FE_PHN562_gl_ram_ram_3_0);
  FE_PHC561_gl_ram_ram_1_0 : CKBD2BWP7T port map(I => FE_PHN489_gl_ram_ram_1_0, Z => FE_PHN561_gl_ram_ram_1_0);
  FE_PHC560_gl_ram_ram_0_1 : CKBD2BWP7T port map(I => FE_PHN506_gl_ram_ram_0_1, Z => FE_PHN560_gl_ram_ram_0_1);
  FE_PHC559_gl_ram_ram_43_0 : BUFFD2BWP7T port map(I => FE_PHN494_gl_ram_ram_43_0, Z => FE_PHN559_gl_ram_ram_43_0);
  FE_PHC558_gl_ram_ram_19_0 : CKBD2BWP7T port map(I => FE_PHN538_gl_ram_ram_19_0, Z => FE_PHN558_gl_ram_ram_19_0);
  FE_PHC557_gl_ram_ram_24_1 : CKBD2BWP7T port map(I => FE_PHN486_gl_ram_ram_24_1, Z => FE_PHN557_gl_ram_ram_24_1);
  FE_PHC556_gl_ram_ram_32_0 : CKBD2BWP7T port map(I => FE_PHN483_gl_ram_ram_32_0, Z => FE_PHN556_gl_ram_ram_32_0);
  FE_PHC555_gl_ram_ram_27_1 : CKBD2BWP7T port map(I => FE_PHN478_gl_ram_ram_27_1, Z => FE_PHN555_gl_ram_ram_27_1);
  FE_PHC554_gl_ram_ram_40_0 : CKBD2BWP7T port map(I => FE_PHN484_gl_ram_ram_40_0, Z => FE_PHN554_gl_ram_ram_40_0);
  FE_PHC553_gl_ram_ram_0_0 : CKBD2BWP7T port map(I => FE_PHN481_gl_ram_ram_0_0, Z => FE_PHN553_gl_ram_ram_0_0);
  FE_PHC552_ml_ms_sr_new_new_data_6 : CKBD0BWP7T port map(I => FE_PHN552_ml_ms_sr_new_new_data_6, Z => FE_PHN468_ml_ms_sr_new_new_data_6);
  FE_PHC551_ml_ms_ed_n_8 : BUFFD3BWP7T port map(I => ml_ms_ed_n_8, Z => FE_PHN551_ml_ms_ed_n_8);
  FE_PHC550_ml_ms_n_34 : CKBD0BWP7T port map(I => ml_ms_n_34, Z => FE_PHN550_ml_ms_n_34);
  FE_PHC549_ml_ms_n_32 : CKBD0BWP7T port map(I => ml_ms_n_32, Z => FE_PHN549_ml_ms_n_32);
  FE_PHC548_ml_ms_n_30 : CKBD0BWP7T port map(I => ml_ms_n_30, Z => FE_PHN548_ml_ms_n_30);
  FE_PHC547_ml_ms_ed_n_5 : DEL02BWP7T port map(I => ml_ms_ed_n_5, Z => FE_PHN547_ml_ms_ed_n_5);
  FE_PHC546_ml_ms_n_58 : DEL01BWP7T port map(I => ml_ms_n_58, Z => FE_PHN546_ml_ms_n_58);
  FE_PHC545_ml_ms_n_21 : CKBD0BWP7T port map(I => FE_PHN545_ml_ms_n_21, Z => ml_ms_n_21);
  FE_PHC544_ml_ms_n_60 : CKBD0BWP7T port map(I => FE_PHN458_ml_ms_n_60, Z => FE_PHN544_ml_ms_n_60);
  FE_PHC543_gl_vgd_horizontal_counter_6 : DEL01BWP7T port map(I => FE_PHN543_gl_vgd_horizontal_counter_6, Z => FE_PHN453_gl_vgd_horizontal_counter_6);
  FE_PHC542_ml_ms_data_sr_11bit_3 : DEL01BWP7T port map(I => FE_PHN542_ml_ms_data_sr_11bit_3, Z => FE_PHN432_ml_ms_data_sr_11bit_3);
  FE_PHC541_gl_ram_ram_8_2 : CKBD0BWP7T port map(I => FE_PHN646_gl_ram_ram_8_2, Z => FE_PHN541_gl_ram_ram_8_2);
  FE_PHC540_gl_ram_ram_25_0 : CKBD0BWP7T port map(I => gl_ram_ram_25(0), Z => FE_PHN540_gl_ram_ram_25_0);
  FE_PHC539_gl_ram_ram_57_1 : CKBD0BWP7T port map(I => gl_ram_ram_57(1), Z => FE_PHN539_gl_ram_ram_57_1);
  FE_PHC538_gl_ram_ram_19_0 : CKBD0BWP7T port map(I => gl_ram_ram_19(0), Z => FE_PHN538_gl_ram_ram_19_0);
  FE_PHC537_gl_ram_ram_50_2 : CKBD0BWP7T port map(I => gl_ram_ram_50(2), Z => FE_PHN537_gl_ram_ram_50_2);
  FE_PHC536_gl_ram_ram_41_0 : CKBD0BWP7T port map(I => FE_PHN626_gl_ram_ram_41_0, Z => FE_PHN536_gl_ram_ram_41_0);
  FE_PHC535_gl_ram_ram_12_2 : CKBD0BWP7T port map(I => gl_ram_ram_12(2), Z => FE_PHN535_gl_ram_ram_12_2);
  FE_PHC534_gl_ram_ram_8_1 : CKBD0BWP7T port map(I => gl_ram_ram_8(1), Z => FE_PHN534_gl_ram_ram_8_1);
  FE_PHC533_gl_ram_ram_48_2 : BUFFD0BWP7T port map(I => gl_ram_ram_48(2), Z => FE_PHN533_gl_ram_ram_48_2);
  FE_PHC532_gl_ram_ram_11_0 : CKBD0BWP7T port map(I => gl_ram_ram_11(0), Z => FE_PHN532_gl_ram_ram_11_0);
  FE_PHC531_gl_ram_ram_89_0 : CKBD0BWP7T port map(I => gl_ram_ram_89(0), Z => FE_PHN531_gl_ram_ram_89_0);
  FE_PHC530_gl_ram_ram_27_0 : CKBD0BWP7T port map(I => FE_PHN639_gl_ram_ram_27_0, Z => FE_PHN530_gl_ram_ram_27_0);
  FE_PHC529_gl_vgd_horizontal_counter_7 : DEL0BWP7T port map(I => gl_vgd_horizontal_counter(7), Z => FE_PHN529_gl_vgd_horizontal_counter_7);
  FE_PHC528_gl_ram_ram_9_2 : BUFFD3BWP7T port map(I => gl_ram_ram_9(2), Z => FE_PHN528_gl_ram_ram_9_2);
  FE_PHC527_gl_ram_ram_40_1 : BUFFD3BWP7T port map(I => gl_ram_ram_40(1), Z => FE_PHN527_gl_ram_ram_40_1);
  FE_PHC526_ml_ms_muxFSM : DEL015BWP7T port map(I => ml_ms_muxFSM, Z => FE_PHN526_ml_ms_muxFSM);
  FE_PHC525_gl_ram_ram_43_1 : BUFFD3BWP7T port map(I => FE_PHN658_gl_ram_ram_43_1, Z => FE_PHN525_gl_ram_ram_43_1);
  FE_PHC524_gl_vgd_horizontal_counter_8 : DEL0BWP7T port map(I => gl_vgd_horizontal_counter(8), Z => FE_PHN524_gl_vgd_horizontal_counter_8);
  FE_PHC523_gl_ram_ram_0_2 : BUFFD3BWP7T port map(I => gl_ram_ram_0(2), Z => FE_PHN523_gl_ram_ram_0_2);
  FE_PHC522_gl_ram_ram_21_0 : CKBD2BWP7T port map(I => gl_ram_ram_21(0), Z => FE_PHN522_gl_ram_ram_21_0);
  FE_PHC521_gl_ram_ram_24_2 : CKBD2BWP7T port map(I => gl_ram_ram_24(2), Z => FE_PHN521_gl_ram_ram_24_2);
  FE_PHC520_gl_ram_ram_58_1 : CKBD2BWP7T port map(I => gl_ram_ram_58(1), Z => FE_PHN520_gl_ram_ram_58_1);
  FE_PHC519_gl_ram_ram_1_2 : CKBD2BWP7T port map(I => gl_ram_ram_1(2), Z => FE_PHN519_gl_ram_ram_1_2);
  FE_PHC518_gl_ram_ram_27_2 : CKBD2BWP7T port map(I => gl_ram_ram_27(2), Z => FE_PHN518_gl_ram_ram_27_2);
  FE_PHC517_gl_ram_ram_2_2 : CKBD2BWP7T port map(I => gl_ram_ram_2(2), Z => FE_PHN517_gl_ram_ram_2_2);
  FE_PHC516_ml_ms_sr_new_new_data_5 : DEL02BWP7T port map(I => ml_ms_sr_new_new_data(5), Z => FE_PHN516_ml_ms_sr_new_new_data_5);
  FE_PHC515_ml_ms_sfsm_state_0 : CKBD0BWP7T port map(I => ml_ms_sfsm_state(0), Z => FE_PHN515_ml_ms_sfsm_state_0);
  FE_PHC514_gl_ram_ram_88_0 : CKBD2BWP7T port map(I => FE_PHN643_gl_ram_ram_88_0, Z => FE_PHN514_gl_ram_ram_88_0);
  FE_PHC513_ml_ms_count_debounce_6 : DEL02BWP7T port map(I => FE_PHN616_ml_ms_count_debounce_6, Z => FE_PHN513_ml_ms_count_debounce_6);
  FE_PHC512_gl_ram_ram_43_2 : DEL02BWP7T port map(I => gl_ram_ram_43(2), Z => FE_PHN512_gl_ram_ram_43_2);
  FE_PHC511_gl_ram_ram_17_1 : DEL02BWP7T port map(I => FE_PHN609_gl_ram_ram_17_1, Z => FE_PHN511_gl_ram_ram_17_1);
  FE_PHC510_gl_ram_ram_11_2 : BUFFD0BWP7T port map(I => FE_PHN573_gl_ram_ram_11_2, Z => FE_PHN510_gl_ram_ram_11_2);
  FE_PHC509_gl_ram_ram_37_2 : BUFFD0BWP7T port map(I => gl_ram_ram_37(2), Z => FE_PHN509_gl_ram_ram_37_2);
  FE_PHC508_gl_ram_ram_11_1 : BUFFD0BWP7T port map(I => gl_ram_ram_11(1), Z => FE_PHN508_gl_ram_ram_11_1);
  FE_PHC507_gl_ram_ram_4_0 : BUFFD0BWP7T port map(I => FE_PHN625_gl_ram_ram_4_0, Z => FE_PHN507_gl_ram_ram_4_0);
  FE_PHC506_gl_ram_ram_0_1 : BUFFD0BWP7T port map(I => gl_ram_ram_0(1), Z => FE_PHN506_gl_ram_ram_0_1);
  FE_PHC505_gl_ram_ram_2_0 : BUFFD0BWP7T port map(I => gl_ram_ram_2(0), Z => FE_PHN505_gl_ram_ram_2_0);
  FE_PHC504_gl_ram_ram_12_1 : BUFFD0BWP7T port map(I => gl_ram_ram_12(1), Z => FE_PHN504_gl_ram_ram_12_1);
  FE_PHC503_gl_ram_ram_3_2 : BUFFD0BWP7T port map(I => gl_ram_ram_3(2), Z => FE_PHN503_gl_ram_ram_3_2);
  FE_PHC502_gl_ram_ram_51_2 : BUFFD0BWP7T port map(I => FE_PHN645_gl_ram_ram_51_2, Z => FE_PHN502_gl_ram_ram_51_2);
  FE_PHC501_gl_ram_ram_56_1 : BUFFD0BWP7T port map(I => gl_ram_ram_56(1), Z => FE_PHN501_gl_ram_ram_56_1);
  FE_PHC500_gl_ram_ram_56_2 : BUFFD0BWP7T port map(I => gl_ram_ram_56(2), Z => FE_PHN500_gl_ram_ram_56_2);
  FE_PHC499_gl_ram_ram_8_0 : CKBD0BWP7T port map(I => gl_ram_ram_8(0), Z => FE_PHN499_gl_ram_ram_8_0);
  FE_PHC498_gl_ram_ram_75_0 : CKBD0BWP7T port map(I => gl_ram_ram_75(0), Z => FE_PHN498_gl_ram_ram_75_0);
  FE_PHC497_gl_ram_ram_32_1 : CKBD0BWP7T port map(I => gl_ram_ram_32(1), Z => FE_PHN497_gl_ram_ram_32_1);
  FE_PHC496_gl_ram_ram_24_0 : BUFFD0BWP7T port map(I => gl_ram_ram_24(0), Z => FE_PHN496_gl_ram_ram_24_0);
  FE_PHC495_gl_ram_ram_29_1 : BUFFD0BWP7T port map(I => gl_ram_ram_29(1), Z => FE_PHN495_gl_ram_ram_29_1);
  FE_PHC494_gl_ram_ram_43_0 : CKBD0BWP7T port map(I => gl_ram_ram_43(0), Z => FE_PHN494_gl_ram_ram_43_0);
  FE_PHC493_gl_ram_ram_35_0 : BUFFD0BWP7T port map(I => gl_ram_ram_35(0), Z => FE_PHN493_gl_ram_ram_35_0);
  FE_PHC492_gl_ram_ram_5_1 : BUFFD0BWP7T port map(I => FE_PHN638_gl_ram_ram_5_1, Z => FE_PHN492_gl_ram_ram_5_1);
  FE_PHC491_gl_ram_ram_9_0 : CKBD0BWP7T port map(I => gl_ram_ram_9(0), Z => FE_PHN491_gl_ram_ram_9_0);
  FE_PHC490_gl_ram_ram_48_1 : BUFFD0BWP7T port map(I => gl_ram_ram_48(1), Z => FE_PHN490_gl_ram_ram_48_1);
  FE_PHC489_gl_ram_ram_1_0 : CKBD0BWP7T port map(I => gl_ram_ram_1(0), Z => FE_PHN489_gl_ram_ram_1_0);
  FE_PHC488_gl_ram_ram_33_0 : BUFFD0BWP7T port map(I => FE_PHN667_gl_ram_ram_33_0, Z => FE_PHN488_gl_ram_ram_33_0);
  FE_PHC487_gl_ram_ram_3_0 : BUFFD0BWP7T port map(I => gl_ram_ram_3(0), Z => FE_PHN487_gl_ram_ram_3_0);
  FE_PHC486_gl_ram_ram_24_1 : CKBD0BWP7T port map(I => gl_ram_ram_24(1), Z => FE_PHN486_gl_ram_ram_24_1);
  FE_PHC485_gl_ram_ram_59_2 : BUFFD0BWP7T port map(I => gl_ram_ram_59(2), Z => FE_PHN485_gl_ram_ram_59_2);
  FE_PHC484_gl_ram_ram_40_0 : BUFFD0BWP7T port map(I => gl_ram_ram_40(0), Z => FE_PHN484_gl_ram_ram_40_0);
  FE_PHC483_gl_ram_ram_32_0 : CKBD0BWP7T port map(I => gl_ram_ram_32(0), Z => FE_PHN483_gl_ram_ram_32_0);
  FE_PHC482_gl_ram_ram_33_2 : CKBD0BWP7T port map(I => FE_PHN631_gl_ram_ram_33_2, Z => FE_PHN482_gl_ram_ram_33_2);
  FE_PHC481_gl_ram_ram_0_0 : CKBD0BWP7T port map(I => gl_ram_ram_0(0), Z => FE_PHN481_gl_ram_ram_0_0);
  FE_PHC480_gl_ram_ram_97_1 : DEL02BWP7T port map(I => gl_ram_ram_97(1), Z => FE_PHN480_gl_ram_ram_97_1);
  FE_PHC479_gl_ram_ram_91_1 : CKBD0BWP7T port map(I => FE_PHN640_gl_ram_ram_91_1, Z => FE_PHN479_gl_ram_ram_91_1);
  FE_PHC478_gl_ram_ram_27_1 : CKBD0BWP7T port map(I => gl_ram_ram_27(1), Z => FE_PHN478_gl_ram_ram_27_1);
  FE_PHC477_gl_ram_ram_35_2 : BUFFD0BWP7T port map(I => gl_ram_ram_35(2), Z => FE_PHN477_gl_ram_ram_35_2);
  FE_PHC476_gl_ram_ram_19_1 : CKBD0BWP7T port map(I => gl_ram_ram_19(1), Z => FE_PHN476_gl_ram_ram_19_1);
  FE_PHC475_gl_ram_ram_34_1 : BUFFD0BWP7T port map(I => FE_PHN649_gl_ram_ram_34_1, Z => FE_PHN475_gl_ram_ram_34_1);
  FE_PHC474_gl_ram_ram_50_1 : CKBD0BWP7T port map(I => gl_ram_ram_50(1), Z => FE_PHN474_gl_ram_ram_50_1);
  FE_PHC473_ml_ms_count_debounce_7 : DEL02BWP7T port map(I => FE_PHN655_ml_ms_count_debounce_7, Z => FE_PHN473_ml_ms_count_debounce_7);
  FE_PHC472_gl_ram_ram_73_2 : BUFFD0BWP7T port map(I => gl_ram_ram_73(2), Z => FE_PHN472_gl_ram_ram_73_2);
  FE_PHC471_gl_ram_n_396 : CKBD0BWP7T port map(I => gl_ram_n_396, Z => FE_PHN471_gl_ram_n_396);
  FE_PHC470_ml_ms_ed_n_2 : CKBD0BWP7T port map(I => ml_ms_ed_n_2, Z => FE_PHN470_ml_ms_ed_n_2);
  FE_PHC469_gl_ram_n_400 : CKBD0BWP7T port map(I => gl_ram_n_400, Z => FE_PHN469_gl_ram_n_400);
  FE_PHC468_ml_ms_sr_new_new_data_6 : DEL02BWP7T port map(I => FE_PHN468_ml_ms_sr_new_new_data_6, Z => ml_ms_sr_new_new_data(6));
  FE_PHC467_ml_ms_mfsm_n_21 : DEL01BWP7T port map(I => ml_ms_mfsm_n_21, Z => FE_PHN467_ml_ms_mfsm_n_21);
  FE_PHC466_ml_ms_sr_new_new_data_7 : DEL02BWP7T port map(I => ml_ms_sr_new_new_data(7), Z => FE_PHN466_ml_ms_sr_new_new_data_7);
  FE_PHC465_gl_gr_lg_local_y_0 : CKBD3BWP7T port map(I => gl_gr_lg_local_y(0), Z => FE_PHN465_gl_gr_lg_local_y_0);
  FE_PHC464_sig_logic_y_0 : DEL01BWP7T port map(I => FE_PHN436_sig_logic_y_0, Z => FE_PHN464_sig_logic_y_0);
  FE_PHC463_ml_ms_count_debounce_10 : CKBD0BWP7T port map(I => FE_PHN433_ml_ms_count_debounce_10, Z => FE_PHN463_ml_ms_count_debounce_10);
  FE_PHC462_gl_ram_ram_82_0 : CKBD0BWP7T port map(I => FE_PHN451_gl_ram_ram_82_0, Z => FE_PHN462_gl_ram_ram_82_0);
  FE_PHC461_ml_il_color1_n_15 : DEL01BWP7T port map(I => FE_PHN437_ml_il_color1_n_15, Z => FE_PHN461_ml_il_color1_n_15);
  FE_PHC460_ml_ms_n_31 : CKBD0BWP7T port map(I => ml_ms_n_31, Z => FE_PHN460_ml_ms_n_31);
  FE_PHC459_ml_ms_n_24 : BUFFD3BWP7T port map(I => ml_ms_n_24, Z => FE_PHN459_ml_ms_n_24);
  FE_PHC458_ml_ms_n_60 : CKBD0BWP7T port map(I => ml_ms_n_60, Z => FE_PHN458_ml_ms_n_60);
  FE_PHC457_ml_ms_n_58 : CKBD0BWP7T port map(I => FE_PHN457_ml_ms_n_58, Z => ml_ms_n_58);
  FE_PHC456_ml_ms_mfsm_n_52 : CKBD0BWP7T port map(I => ml_ms_mfsm_n_52, Z => FE_PHN456_ml_ms_mfsm_n_52);
  FE_PHC455_gl_gr_lg_lv_n_15 : DEL0BWP7T port map(I => gl_gr_lg_lv_n_15, Z => FE_PHN455_gl_gr_lg_lv_n_15);
  FE_PHC454_ml_ms_mfsm_n_0 : DEL01BWP7T port map(I => ml_ms_mfsm_n_0, Z => FE_PHN454_ml_ms_mfsm_n_0);
  FE_PHC453_gl_vgd_horizontal_counter_6 : DEL0BWP7T port map(I => FE_PHN453_gl_vgd_horizontal_counter_6, Z => gl_vgd_horizontal_counter(6));
  FE_PHC452_ml_ms_count25M_8 : DEL01BWP7T port map(I => FE_PHN452_ml_ms_count25M_8, Z => FE_PHN332_ml_ms_count25M_8);
  FE_PHC451_gl_ram_ram_82_0 : CKBD0BWP7T port map(I => gl_ram_ram_82(0), Z => FE_PHN451_gl_ram_ram_82_0);
  FE_PHC450_gl_ram_ram_20_2 : DEL01BWP7T port map(I => FE_PHN310_gl_ram_ram_20_2, Z => FE_PHN450_gl_ram_ram_20_2);
  FE_PHC449_gl_ram_ram_46_2 : DEL01BWP7T port map(I => FE_PHN314_gl_ram_ram_46_2, Z => FE_PHN449_gl_ram_ram_46_2);
  FE_PHC448_ml_ms_tb_n_0 : DEL01BWP7T port map(I => FE_PHN448_ml_ms_tb_n_0, Z => ml_ms_tb_n_0);
  FE_PHC447_gl_ram_ram_37_0 : DEL01BWP7T port map(I => gl_ram_ram_37(0), Z => FE_PHN447_gl_ram_ram_37_0);
  FE_PHC446_ml_ms_mux_select : DEL02BWP7T port map(I => ml_ms_mux_select, Z => FE_PHN446_ml_ms_mux_select);
  FE_PHC445_gl_gr_lg_lcountdown_n_2 : DEL01BWP7T port map(I => FE_PHN445_gl_gr_lg_lcountdown_n_2, Z => gl_gr_lg_lcountdown_n_2);
  FE_PHC444_gl_ram_ram_80_0 : DEL01BWP7T port map(I => FE_PHN312_gl_ram_ram_80_0, Z => FE_PHN444_gl_ram_ram_80_0);
  FE_PHC443_gl_gr_lg_lcountdown_n_4 : DEL01BWP7T port map(I => gl_gr_lg_lcountdown_n_4, Z => FE_PHN443_gl_gr_lg_lcountdown_n_4);
  FE_PHC442_gl_ram_ram_5_0 : DEL01BWP7T port map(I => FE_PHN311_gl_ram_ram_5_0, Z => FE_PHN442_gl_ram_ram_5_0);
  FE_PHC441_ml_ms_n_2 : DEL02BWP7T port map(I => ml_ms_n_2, Z => FE_PHN441_ml_ms_n_2);
  FE_PHC440_gl_ram_ram_86_1 : DEL01BWP7T port map(I => gl_ram_ram_86(1), Z => FE_PHN440_gl_ram_ram_86_1);
  FE_PHC439_gl_ram_ram_61_1 : DEL01BWP7T port map(I => FE_PHN315_gl_ram_ram_61_1, Z => FE_PHN439_gl_ram_ram_61_1);
  FE_PHC438_gl_ram_ram_10_0 : DEL01BWP7T port map(I => FE_PHN316_gl_ram_ram_10_0, Z => FE_PHN438_gl_ram_ram_10_0);
  FE_PHC437_ml_il_color1_n_15 : CKBD0BWP7T port map(I => ml_il_color1_n_15, Z => FE_PHN437_ml_il_color1_n_15);
  FE_PHC436_sig_logic_y_0 : CKBD0BWP7T port map(I => sig_logic_y(0), Z => FE_PHN436_sig_logic_y_0);
  FE_PHC435_gl_gr_lg_lcountdown_n_15 : BUFFD5BWP7T port map(I => gl_gr_lg_lcountdown_n_15, Z => FE_PHN435_gl_gr_lg_lcountdown_n_15);
  FE_PHC434_ml_ms_count_debounce_6 : DEL02BWP7T port map(I => FE_PHN434_ml_ms_count_debounce_6, Z => ml_ms_count_debounce(6));
  FE_PHC433_ml_ms_count_debounce_10 : DEL02BWP7T port map(I => ml_ms_count_debounce(10), Z => FE_PHN433_ml_ms_count_debounce_10);
  FE_PHC432_ml_ms_data_sr_11bit_3 : CKBD0BWP7T port map(I => FE_PHN432_ml_ms_data_sr_11bit_3, Z => FE_PHN275_ml_ms_data_sr_11bit_3);
  FE_PHC431_gl_ram_ram_60_0 : DEL0BWP7T port map(I => gl_ram_ram_60(0), Z => FE_PHN431_gl_ram_ram_60_0);
  FE_PHC430_gl_ram_ram_60_2 : DEL0BWP7T port map(I => gl_ram_ram_60(2), Z => FE_PHN430_gl_ram_ram_60_2);
  FE_PHC429_gl_ram_ram_60_1 : DEL0BWP7T port map(I => gl_ram_ram_60(1), Z => FE_PHN429_gl_ram_ram_60_1);
  FE_PHC428_gl_ram_ram_36_2 : DEL0BWP7T port map(I => gl_ram_ram_36(2), Z => FE_PHN428_gl_ram_ram_36_2);
  FE_PHC427_gl_ram_ram_33_1 : DEL0BWP7T port map(I => gl_ram_ram_33(1), Z => FE_PHN427_gl_ram_ram_33_1);
  FE_PHC426_gl_ram_ram_96_2 : DEL0BWP7T port map(I => gl_ram_ram_96(2), Z => FE_PHN426_gl_ram_ram_96_2);
  FE_PHC425_gl_ram_n_495 : DEL0BWP7T port map(I => gl_ram_n_495, Z => FE_PHN425_gl_ram_n_495);
  FE_PHC424_gl_ram_ram_31_2 : DEL0BWP7T port map(I => gl_ram_ram_31(2), Z => FE_PHN424_gl_ram_ram_31_2);
  FE_PHC423_gl_ram_ram_25_1 : DEL0BWP7T port map(I => gl_ram_ram_25(1), Z => FE_PHN423_gl_ram_ram_25_1);
  FE_PHC422_gl_ram_ram_20_1 : DEL0BWP7T port map(I => gl_ram_ram_20(1), Z => FE_PHN422_gl_ram_ram_20_1);
  FE_PHC421_gl_ram_ram_65_2 : DEL0BWP7T port map(I => gl_ram_ram_65(2), Z => FE_PHN421_gl_ram_ram_65_2);
  FE_PHC420_gl_ram_ram_97_0 : DEL0BWP7T port map(I => gl_ram_ram_97(0), Z => FE_PHN420_gl_ram_ram_97_0);
  FE_PHC419_gl_ram_ram_96_1 : DEL0BWP7T port map(I => gl_ram_ram_96(1), Z => FE_PHN419_gl_ram_ram_96_1);
  FE_PHC418_gl_ram_ram_83_0 : DEL0BWP7T port map(I => gl_ram_ram_83(0), Z => FE_PHN418_gl_ram_ram_83_0);
  FE_PHC417_gl_ram_ram_73_0 : DEL0BWP7T port map(I => gl_ram_ram_73(0), Z => FE_PHN417_gl_ram_ram_73_0);
  FE_PHC416_gl_ram_ram_66_0 : DEL0BWP7T port map(I => gl_ram_ram_66(0), Z => FE_PHN416_gl_ram_ram_66_0);
  FE_PHC415_gl_ram_n_496 : DEL0BWP7T port map(I => gl_ram_n_496, Z => FE_PHN415_gl_ram_n_496);
  FE_PHC414_gl_ram_ram_67_0 : DEL0BWP7T port map(I => gl_ram_ram_67(0), Z => FE_PHN414_gl_ram_ram_67_0);
  FE_PHC413_gl_ram_n_394 : DEL0BWP7T port map(I => gl_ram_n_394, Z => FE_PHN413_gl_ram_n_394);
  FE_PHC412_gl_ram_ram_73_1 : DEL0BWP7T port map(I => gl_ram_ram_73(1), Z => FE_PHN412_gl_ram_ram_73_1);
  FE_PHC411_gl_ram_ram_41_2 : DEL0BWP7T port map(I => gl_ram_ram_41(2), Z => FE_PHN411_gl_ram_ram_41_2);
  FE_PHC410_ml_ms_cnt_count_0 : DEL0BWP7T port map(I => ml_ms_cnt_count(0), Z => FE_PHN410_ml_ms_cnt_count_0);
  FE_PHC409_gl_ram_ram_98_2 : DEL0BWP7T port map(I => gl_ram_ram_98(2), Z => FE_PHN409_gl_ram_ram_98_2);
  FE_PHC408_gl_ram_ram_82_1 : DEL0BWP7T port map(I => gl_ram_ram_82(1), Z => FE_PHN408_gl_ram_ram_82_1);
  FE_PHC407_gl_gr_lg_lv_n_3 : DEL0BWP7T port map(I => gl_gr_lg_lv_n_3, Z => FE_PHN407_gl_gr_lg_lv_n_3);
  FE_PHC406_ml_il_color1_state_hs_1 : DEL0BWP7T port map(I => FE_PHN406_ml_il_color1_state_hs_1, Z => ml_il_color1_state_hs(1));
  FE_PHC405_gl_gr_lg_lcountdown_n_13 : DEL0BWP7T port map(I => gl_gr_lg_lcountdown_n_13, Z => FE_PHN405_gl_gr_lg_lcountdown_n_13);
  FE_PHC404_gl_gr_lg_lcountdown_n_17 : DEL0BWP7T port map(I => gl_gr_lg_lcountdown_n_17, Z => FE_PHN404_gl_gr_lg_lcountdown_n_17);
  FE_PHC403_gl_gr_lg_lcountdown_n_19 : DEL0BWP7T port map(I => gl_gr_lg_lcountdown_n_19, Z => FE_PHN403_gl_gr_lg_lcountdown_n_19);
  FE_PHC402_gl_gr_lg_lcountdown_n_8 : DEL0BWP7T port map(I => gl_gr_lg_lcountdown_n_8, Z => FE_PHN402_gl_gr_lg_lcountdown_n_8);
  FE_PHC401_gl_gr_lg_lcountdown_n_20 : DEL0BWP7T port map(I => gl_gr_lg_lcountdown_n_20, Z => FE_PHN401_gl_gr_lg_lcountdown_n_20);
  FE_PHC400_gl_gr_lg_lcountdown_n_11 : DEL0BWP7T port map(I => FE_PHN400_gl_gr_lg_lcountdown_n_11, Z => gl_gr_lg_lcountdown_n_11);
  FE_PHC399_gl_gr_lg_lcountdown_n_21 : DEL0BWP7T port map(I => gl_gr_lg_lcountdown_n_21, Z => FE_PHN399_gl_gr_lg_lcountdown_n_21);
  FE_PHC398_gl_gr_lg_lcountdown_n_0 : DEL0BWP7T port map(I => gl_gr_lg_lcountdown_n_0, Z => FE_PHN398_gl_gr_lg_lcountdown_n_0);
  FE_PHC397_ml_ms_cntD_n_19 : DEL0BWP7T port map(I => ml_ms_cntD_n_19, Z => FE_PHN397_ml_ms_cntD_n_19);
  FE_PHC396_gl_gr_lg_lcountdown_sig_edge_fall : DEL02BWP7T port map(I => gl_gr_lg_lcountdown_sig_edge_fall, Z => FE_PHN396_gl_gr_lg_lcountdown_sig_edge_fall);
  FE_PHC395_ml_il_x1_n_9 : DEL02BWP7T port map(I => ml_il_x1_n_9, Z => FE_PHN395_ml_il_x1_n_9);
  FE_PHC394_ml_ms_mfsm_n_44 : DEL0BWP7T port map(I => ml_ms_mfsm_n_44, Z => FE_PHN394_ml_ms_mfsm_n_44);
  FE_PHC393_ml_ms_cnt_n_5 : DEL0BWP7T port map(I => ml_ms_cnt_n_5, Z => FE_PHN393_ml_ms_cnt_n_5);
  FE_PHC392_gl_ram_n_145 : DEL0BWP7T port map(I => gl_ram_n_145, Z => FE_PHN392_gl_ram_n_145);
  FE_PHC391_ml_ms_tb_n_5 : DEL0BWP7T port map(I => FE_PHN391_ml_ms_tb_n_5, Z => ml_ms_tb_n_5);
  FE_PHC390_ml_ms_cnt_n_9 : DEL0BWP7T port map(I => ml_ms_cnt_n_9, Z => FE_PHN390_ml_ms_cnt_n_9);
  FE_PHC389_gl_ram_n_563 : DEL0BWP7T port map(I => gl_ram_n_563, Z => FE_PHN389_gl_ram_n_563);
  FE_PHC388_ml_ms_tb_n_6 : DEL0BWP7T port map(I => FE_PHN388_ml_ms_tb_n_6, Z => ml_ms_tb_n_6);
  FE_PHC387_ml_ms_mfsm_n_38 : DEL0BWP7T port map(I => ml_ms_mfsm_n_38, Z => FE_PHN387_ml_ms_mfsm_n_38);
  FE_PHC386_ml_ms_cnt_n_7 : DEL0BWP7T port map(I => ml_ms_cnt_n_7, Z => FE_PHN386_ml_ms_cnt_n_7);
  FE_PHC385_ml_il_color1_n_14 : DEL0BWP7T port map(I => FE_PHN385_ml_il_color1_n_14, Z => ml_il_color1_n_14);
  FE_PHC384_ml_il_y1_n_9 : DEL02BWP7T port map(I => ml_il_y1_n_9, Z => FE_PHN384_ml_il_y1_n_9);
  FE_PHC383_ml_ms_cnt_n_3 : DEL0BWP7T port map(I => ml_ms_cnt_n_3, Z => FE_PHN383_ml_ms_cnt_n_3);
  FE_PHC382_gl_ram_n_564 : DEL0BWP7T port map(I => gl_ram_n_564, Z => FE_PHN382_gl_ram_n_564);
  FE_PHC381_gl_ram_n_567 : DEL1BWP7T port map(I => FE_PHN381_gl_ram_n_567, Z => gl_ram_n_567);
  FE_PHC380_gl_gr_lg_lv_n_12 : DEL0BWP7T port map(I => gl_gr_lg_lv_n_12, Z => FE_PHN380_gl_gr_lg_lv_n_12);
  FE_PHC379_ml_ms_n_54 : DEL0BWP7T port map(I => FE_PHN379_ml_ms_n_54, Z => ml_ms_n_54);
  FE_PHC378_ml_il_color1_n_13 : DEL0BWP7T port map(I => ml_il_color1_n_13, Z => FE_PHN378_ml_il_color1_n_13);
  FE_PHC377_gl_ram_n_247 : DEL1BWP7T port map(I => gl_ram_n_247, Z => FE_PHN377_gl_ram_n_247);
  FE_PHC376_gl_ram_n_308 : DEL1BWP7T port map(I => gl_ram_n_308, Z => FE_PHN376_gl_ram_n_308);
  FE_PHC375_gl_ram_n_552 : DEL0BWP7T port map(I => gl_ram_n_552, Z => FE_PHN375_gl_ram_n_552);
  FE_PHC374_ml_il_color1_n_10 : DEL0BWP7T port map(I => FE_PHN374_ml_il_color1_n_10, Z => ml_il_color1_n_10);
  FE_PHC373_ml_ms_cnt_n_21 : DEL0BWP7T port map(I => ml_ms_cnt_n_21, Z => FE_PHN373_ml_ms_cnt_n_21);
  FE_PHC372_ml_ms_n_57 : DEL0BWP7T port map(I => ml_ms_n_57, Z => FE_PHN372_ml_ms_n_57);
  FE_PHC371_gl_vgd_n_64 : DEL1BWP7T port map(I => gl_vgd_n_64, Z => FE_PHN371_gl_vgd_n_64);
  FE_PHC370_gl_ram_n_243 : DEL1BWP7T port map(I => gl_ram_n_243, Z => FE_PHN370_gl_ram_n_243);
  FE_PHC369_gl_ram_n_237 : DEL0BWP7T port map(I => gl_ram_n_237, Z => FE_PHN369_gl_ram_n_237);
  FE_PHC368_ml_ms_cnt_n_22 : DEL0BWP7T port map(I => ml_ms_cnt_n_22, Z => FE_PHN368_ml_ms_cnt_n_22);
  FE_PHC367_ml_ms_mfsm_n_36 : DEL0BWP7T port map(I => ml_ms_mfsm_n_36, Z => FE_PHN367_ml_ms_mfsm_n_36);
  FE_PHC366_gl_ram_n_568 : DEL0BWP7T port map(I => gl_ram_n_568, Z => FE_PHN366_gl_ram_n_568);
  FE_PHC365_gl_ram_n_80 : DEL1BWP7T port map(I => FE_PHN365_gl_ram_n_80, Z => gl_ram_n_80);
  FE_PHC364_gl_gr_lg_lv_n_14 : DEL1BWP7T port map(I => gl_gr_lg_lv_n_14, Z => FE_PHN364_gl_gr_lg_lv_n_14);
  FE_PHC363_ml_ms_cnt_n_19 : DEL0BWP7T port map(I => FE_PHN363_ml_ms_cnt_n_19, Z => ml_ms_cnt_n_19);
  FE_PHC362_gl_sig_v : DEL1BWP7T port map(I => gl_sig_v, Z => FE_PHN362_gl_sig_v);
  FE_PHC361_gl_ram_n_78 : DEL1BWP7T port map(I => gl_ram_n_78, Z => FE_PHN361_gl_ram_n_78);
  FE_PHC360_gl_ram_n_142 : DEL1BWP7T port map(I => gl_ram_n_142, Z => FE_PHN360_gl_ram_n_142);
  FE_PHC359_gl_ram_n_77 : DEL1BWP7T port map(I => gl_ram_n_77, Z => FE_PHN359_gl_ram_n_77);
  FE_PHC358_gl_sig_scale_v : DEL1BWP7T port map(I => FE_PHN358_gl_sig_scale_v, Z => gl_sig_scale_v);
  FE_PHC357_gl_sig_scale_h : DEL1BWP7T port map(I => gl_sig_scale_h, Z => FE_PHN357_gl_sig_scale_h);
  FE_PHC356_gl_gr_lg_sig_countdown_10 : DEL02BWP7T port map(I => FE_PHN356_gl_gr_lg_sig_countdown_10, Z => gl_gr_lg_sig_countdown(10));
  FE_PHC355_gl_gr_lg_sig_countdown_5 : DEL02BWP7T port map(I => gl_gr_lg_sig_countdown(5), Z => FE_PHN355_gl_gr_lg_sig_countdown_5);
  FE_PHC354_gl_gr_lg_sig_countdown_2 : DEL0BWP7T port map(I => gl_gr_lg_sig_countdown(2), Z => FE_PHN354_gl_gr_lg_sig_countdown_2);
  FE_PHC353_gl_gr_lg_sig_countdown_0 : CKBD0BWP7T port map(I => gl_gr_lg_sig_countdown(0), Z => FE_PHN353_gl_gr_lg_sig_countdown_0);
  FE_PHC352_gl_gr_lg_sig_countdown_1 : DEL02BWP7T port map(I => gl_gr_lg_sig_countdown(1), Z => FE_PHN352_gl_gr_lg_sig_countdown_1);
  FE_PHC351_sig_logic_x_0 : DEL1BWP7T port map(I => FE_PHN351_sig_logic_x_0, Z => sig_logic_x(0));
  FE_PHC350_ml_ms_mfsm_state_4 : DEL02BWP7T port map(I => ml_ms_mfsm_state(4), Z => FE_PHN350_ml_ms_mfsm_state_4);
  FE_PHC349_sig_logic_y_0 : DEL02BWP7T port map(I => FE_PHN349_sig_logic_y_0, Z => sig_logic_y(0));
  FE_PHC348_gl_gr_lg_local_y_0 : DEL02BWP7T port map(I => FE_PHN348_gl_gr_lg_local_y_0, Z => gl_gr_lg_local_y(0));
  FE_PHC347_ml_ms_mfsm_state_3 : CKBD0BWP7T port map(I => ml_ms_mfsm_state(3), Z => FE_PHN347_ml_ms_mfsm_state_3);
  FE_PHC346_gl_vgd_horizontal_counter_4 : DEL1BWP7T port map(I => FE_PHN346_gl_vgd_horizontal_counter_4, Z => gl_vgd_horizontal_counter(4));
  FE_PHC345_gl_vgd_horizontal_counter_1 : DEL1BWP7T port map(I => gl_vgd_horizontal_counter(1), Z => FE_PHN345_gl_vgd_horizontal_counter_1);
  FE_PHC344_gl_vgd_horizontal_counter_2 : DEL1BWP7T port map(I => gl_vgd_horizontal_counter(2), Z => FE_PHN344_gl_vgd_horizontal_counter_2);
  FE_PHC343_gl_vgd_horizontal_counter_5 : DEL1BWP7T port map(I => gl_vgd_horizontal_counter(5), Z => FE_PHN343_gl_vgd_horizontal_counter_5);
  FE_PHC342_gl_vgd_horizontal_counter_3 : DEL1BWP7T port map(I => FE_PHN342_gl_vgd_horizontal_counter_3, Z => gl_vgd_horizontal_counter(3));
  FE_PHC341_ml_ms_cnt_count_1 : DEL0BWP7T port map(I => ml_ms_cnt_count(1), Z => FE_PHN341_ml_ms_cnt_count_1);
  FE_PHC340_gl_vgd_horizontal_counter_0 : DEL1BWP7T port map(I => gl_vgd_horizontal_counter(0), Z => FE_PHN340_gl_vgd_horizontal_counter_0);
  FE_PHC339_gl_vgd_horizontal_counter_9 : DEL1BWP7T port map(I => FE_PHN339_gl_vgd_horizontal_counter_9, Z => gl_vgd_horizontal_counter(9));
  FE_PHC338_ml_ms_mfsm_state_2 : DEL02BWP7T port map(I => ml_ms_mfsm_state(2), Z => FE_PHN338_ml_ms_mfsm_state_2);
  FE_PHC337_gl_vgd_vertical_counter_2 : DEL1BWP7T port map(I => FE_PHN337_gl_vgd_vertical_counter_2, Z => gl_vgd_vertical_counter(2));
  FE_PHC336_gl_vgd_vertical_counter_0 : DEL1BWP7T port map(I => FE_PHN336_gl_vgd_vertical_counter_0, Z => gl_vgd_vertical_counter(0));
  FE_PHC335_ml_ms_count15k_1 : DEL02BWP7T port map(I => ml_ms_count15k(1), Z => FE_PHN335_ml_ms_count15k_1);
  FE_PHC334_ml_ms_count15k_0 : DEL02BWP7T port map(I => FE_PHN334_ml_ms_count15k_0, Z => ml_ms_count15k(0));
  FE_PHC333_gl_vgd_vertical_counter_1 : DEL1BWP7T port map(I => FE_PHN333_gl_vgd_vertical_counter_1, Z => gl_vgd_vertical_counter(1));
  FE_PHC332_ml_ms_count25M_8 : DEL02BWP7T port map(I => FE_PHN332_ml_ms_count25M_8, Z => ml_ms_count25M(8));
  FE_PHC331_gl_vgd_vertical_counter_9 : DEL1BWP7T port map(I => FE_PHN331_gl_vgd_vertical_counter_9, Z => gl_vgd_vertical_counter(9));
  FE_PHC330_gl_vgd_vertical_counter_6 : DEL1BWP7T port map(I => FE_PHN330_gl_vgd_vertical_counter_6, Z => gl_vgd_vertical_counter(6));
  FE_PHC329_ml_ms_mfsm_n_53 : DEL0BWP7T port map(I => ml_ms_mfsm_n_53, Z => FE_PHN329_ml_ms_mfsm_n_53);
  FE_PHC328_gl_vgd_vertical_counter_7 : DEL1BWP7T port map(I => FE_PHN328_gl_vgd_vertical_counter_7, Z => gl_vgd_vertical_counter(7));
  FE_PHC327_gl_ram_n_5 : DEL1BWP7T port map(I => gl_ram_n_5, Z => FE_PHN327_gl_ram_n_5);
  FE_PHC326_gl_vgd_vertical_counter_5 : DEL1BWP7T port map(I => gl_vgd_vertical_counter(5), Z => FE_PHN326_gl_vgd_vertical_counter_5);
  FE_PHC325_gl_gr_lg_lv_sig_edges : DEL0BWP7T port map(I => gl_gr_lg_lv_sig_edges, Z => FE_PHN325_gl_gr_lg_lv_sig_edges);
  FE_PHC324_gl_vgd_vertical_counter_4 : DEL1BWP7T port map(I => gl_vgd_vertical_counter(4), Z => FE_PHN324_gl_vgd_vertical_counter_4);
  FE_PHC323_ml_ms_count25M_9 : DEL0BWP7T port map(I => ml_ms_count25M(9), Z => FE_PHN323_ml_ms_count25M_9);
  FE_PHC322_gl_vgd_vertical_counter_3 : DEL1BWP7T port map(I => FE_PHN322_gl_vgd_vertical_counter_3, Z => gl_vgd_vertical_counter(3));
  FE_PHC321_gl_vgd_n_77 : DEL1BWP7T port map(I => gl_vgd_n_77, Z => FE_PHN321_gl_vgd_n_77);
  FE_PHC320_ml_buttons_mouse_3 : DEL1BWP7T port map(I => ml_buttons_mouse(3), Z => FE_PHN320_ml_buttons_mouse_3);
  FE_PHC319_gl_gr_lg_sig_countdown_3 : DEL02BWP7T port map(I => gl_gr_lg_sig_countdown(3), Z => FE_PHN319_gl_gr_lg_sig_countdown_3);
  FE_PHC318_ml_ms_count25M_6 : DEL0BWP7T port map(I => ml_ms_count25M(6), Z => FE_PHN318_ml_ms_count25M_6);
  FE_PHC317_gl_ram_ram_86_1 : DEL0BWP7T port map(I => FE_PHN440_gl_ram_ram_86_1, Z => FE_PHN317_gl_ram_ram_86_1);
  FE_PHC316_gl_ram_ram_10_0 : DEL0BWP7T port map(I => gl_ram_ram_10(0), Z => FE_PHN316_gl_ram_ram_10_0);
  FE_PHC315_gl_ram_ram_61_1 : DEL0BWP7T port map(I => gl_ram_ram_61(1), Z => FE_PHN315_gl_ram_ram_61_1);
  FE_PHC314_gl_ram_ram_46_2 : DEL0BWP7T port map(I => gl_ram_ram_46(2), Z => FE_PHN314_gl_ram_ram_46_2);
  FE_PHC313_ml_ms_cntD_count_1 : DEL0BWP7T port map(I => FE_PHN313_ml_ms_cntD_count_1, Z => ml_ms_cntD_count(1));
  FE_PHC312_gl_ram_ram_80_0 : DEL0BWP7T port map(I => gl_ram_ram_80(0), Z => FE_PHN312_gl_ram_ram_80_0);
  FE_PHC311_gl_ram_ram_5_0 : DEL0BWP7T port map(I => gl_ram_ram_5(0), Z => FE_PHN311_gl_ram_ram_5_0);
  FE_PHC310_gl_ram_ram_20_2 : DEL0BWP7T port map(I => gl_ram_ram_20(2), Z => FE_PHN310_gl_ram_ram_20_2);
  FE_PHC309_gl_ram_ram_37_0 : DEL0BWP7T port map(I => FE_PHN447_gl_ram_ram_37_0, Z => FE_PHN309_gl_ram_ram_37_0);
  FE_PHC308_ml_ms_count25M_5 : CKBD0BWP7T port map(I => ml_ms_count25M(5), Z => FE_PHN308_ml_ms_count25M_5);
  FE_PHC307_data_in : DEL0BWP7T port map(I => data_in, Z => FE_PHN307_data_in);
  FE_PHC306_gl_ram_ram_39_2 : DEL2BWP7T port map(I => gl_ram_ram_39(2), Z => FE_PHN306_gl_ram_ram_39_2);
  FE_PHC305_gl_ram_ram_70_2 : DEL2BWP7T port map(I => gl_ram_ram_70(2), Z => FE_PHN305_gl_ram_ram_70_2);
  FE_PHC304_gl_gr_lg_lcountdown_l_edge_reg1 : DEL1BWP7T port map(I => gl_gr_lg_lcountdown_l_edge_reg1, Z => FE_PHN304_gl_gr_lg_lcountdown_l_edge_reg1);
  FE_PHC303_gl_ram_ram_71_1 : DEL2BWP7T port map(I => gl_ram_ram_71(1), Z => FE_PHN303_gl_ram_ram_71_1);
  FE_PHC302_gl_ram_ram_87_2 : DEL2BWP7T port map(I => gl_ram_ram_87(2), Z => FE_PHN302_gl_ram_ram_87_2);
  FE_PHC301_gl_gr_lg_lh_n_21 : DEL1BWP7T port map(I => gl_gr_lg_lh_n_21, Z => FE_PHN301_gl_gr_lg_lh_n_21);
  FE_PHC300_gl_gr_lg_lh_n_14 : DEL1BWP7T port map(I => gl_gr_lg_lh_n_14, Z => FE_PHN300_gl_gr_lg_lh_n_14);
  FE_PHC299_ml_ms_data_sr_11bit_7 : DEL0BWP7T port map(I => FE_PHN299_ml_ms_data_sr_11bit_7, Z => ml_ms_data_sr_11bit(7));
  FE_PHC298_gl_ram_ram_86_2 : DEL1BWP7T port map(I => gl_ram_ram_86(2), Z => FE_PHN298_gl_ram_ram_86_2);
  FE_PHC297_gl_Hint : DEL0BWP7T port map(I => FE_PHN297_gl_Hint, Z => gl_Hint);
  FE_PHC296_gl_ram_ram_78_1 : DEL1BWP7T port map(I => gl_ram_ram_78(1), Z => FE_PHN296_gl_ram_ram_78_1);
  FE_PHC295_gl_ram_ram_14_2 : DEL1BWP7T port map(I => gl_ram_ram_14(2), Z => FE_PHN295_gl_ram_ram_14_2);
  FE_PHC294_gl_ram_ram_82_2 : DEL1BWP7T port map(I => gl_ram_ram_82(2), Z => FE_PHN294_gl_ram_ram_82_2);
  FE_PHC293_gl_ram_ram_39_0 : DEL1BWP7T port map(I => gl_ram_ram_39(0), Z => FE_PHN293_gl_ram_ram_39_0);
  FE_PHC292_gl_ram_ram_14_0 : DEL1BWP7T port map(I => gl_ram_ram_14(0), Z => FE_PHN292_gl_ram_ram_14_0);
  FE_PHC291_gl_ram_ram_86_0 : DEL1BWP7T port map(I => gl_ram_ram_86(0), Z => FE_PHN291_gl_ram_ram_86_0);
  FE_PHC290_gl_ram_ram_53_0 : DEL1BWP7T port map(I => gl_ram_ram_53(0), Z => FE_PHN290_gl_ram_ram_53_0);
  FE_PHC289_gl_ram_ram_46_1 : DEL1BWP7T port map(I => gl_ram_ram_46(1), Z => FE_PHN289_gl_ram_ram_46_1);
  FE_PHC288_gl_ram_ram_38_1 : DEL1BWP7T port map(I => gl_ram_ram_38(1), Z => FE_PHN288_gl_ram_ram_38_1);
  FE_PHC287_gl_ram_ram_23_2 : DEL1BWP7T port map(I => gl_ram_ram_23(2), Z => FE_PHN287_gl_ram_ram_23_2);
  FE_PHC286_gl_ram_ram_76_0 : DEL1BWP7T port map(I => gl_ram_ram_76(0), Z => FE_PHN286_gl_ram_ram_76_0);
  FE_PHC285_gl_ram_ram_36_1 : DEL1BWP7T port map(I => gl_ram_ram_36(1), Z => FE_PHN285_gl_ram_ram_36_1);
  FE_PHC284_ml_mouseY_0 : DEL2BWP7T port map(I => ml_mouseY(0), Z => FE_PHN284_ml_mouseY_0);
  FE_PHC283_gl_ram_ram_53_1 : DEL1BWP7T port map(I => gl_ram_ram_53(1), Z => FE_PHN283_gl_ram_ram_53_1);
  FE_PHC282_gl_ram_ram_23_1 : DEL1BWP7T port map(I => gl_ram_ram_23(1), Z => FE_PHN282_gl_ram_ram_23_1);
  FE_PHC281_gl_ram_ram_22_1 : DEL1BWP7T port map(I => gl_ram_ram_22(1), Z => FE_PHN281_gl_ram_ram_22_1);
  FE_PHC280_gl_ram_ram_66_2 : DEL1BWP7T port map(I => gl_ram_ram_66(2), Z => FE_PHN280_gl_ram_ram_66_2);
  FE_PHC279_ml_ms_data_sr_11bit_2 : DEL1BWP7T port map(I => ml_ms_data_sr_11bit(2), Z => FE_PHN279_ml_ms_data_sr_11bit_2);
  FE_PHC278_gl_ram_ram_52_2 : DEL1BWP7T port map(I => gl_ram_ram_52(2), Z => FE_PHN278_gl_ram_ram_52_2);
  FE_PHC277_gl_ram_ram_63_1 : DEL1BWP7T port map(I => gl_ram_ram_63(1), Z => FE_PHN277_gl_ram_ram_63_1);
  FE_PHC276_gl_ram_ram_55_1 : DEL1BWP7T port map(I => gl_ram_ram_55(1), Z => FE_PHN276_gl_ram_ram_55_1);
  FE_PHC275_ml_ms_data_sr_11bit_3 : DEL02BWP7T port map(I => FE_PHN275_ml_ms_data_sr_11bit_3, Z => ml_ms_data_sr_11bit(3));
  FE_PHC274_gl_ram_ram_36_0 : DEL1BWP7T port map(I => gl_ram_ram_36(0), Z => FE_PHN274_gl_ram_ram_36_0);
  FE_PHC273_gl_ram_ram_63_0 : DEL1BWP7T port map(I => gl_ram_ram_63(0), Z => FE_PHN273_gl_ram_ram_63_0);
  FE_PHC272_gl_ram_ram_47_0 : DEL1BWP7T port map(I => gl_ram_ram_47(0), Z => FE_PHN272_gl_ram_ram_47_0);
  FE_PHC271_gl_ram_ram_87_1 : DEL1BWP7T port map(I => gl_ram_ram_87(1), Z => FE_PHN271_gl_ram_ram_87_1);
  FE_PHC270_gl_ram_ram_76_2 : DEL1BWP7T port map(I => gl_ram_ram_76(2), Z => FE_PHN270_gl_ram_ram_76_2);
  FE_PHC269_gl_ram_ram_6_0 : DEL1BWP7T port map(I => gl_ram_ram_6(0), Z => FE_PHN269_gl_ram_ram_6_0);
  FE_PHC268_gl_ram_ram_6_1 : DEL1BWP7T port map(I => gl_ram_ram_6(1), Z => FE_PHN268_gl_ram_ram_6_1);
  FE_PHC267_gl_ram_ram_15_2 : DEL1BWP7T port map(I => gl_ram_ram_15(2), Z => FE_PHN267_gl_ram_ram_15_2);
  FE_PHC266_gl_ram_ram_13_0 : DEL1BWP7T port map(I => gl_ram_ram_13(0), Z => FE_PHN266_gl_ram_ram_13_0);
  FE_PHC265_gl_ram_ram_22_0 : DEL1BWP7T port map(I => gl_ram_ram_22(0), Z => FE_PHN265_gl_ram_ram_22_0);
  FE_PHC264_gl_ram_ram_68_0 : DEL1BWP7T port map(I => gl_ram_ram_68(0), Z => FE_PHN264_gl_ram_ram_68_0);
  FE_PHC263_gl_ram_ram_6_2 : DEL1BWP7T port map(I => gl_ram_ram_6(2), Z => FE_PHN263_gl_ram_ram_6_2);
  FE_PHC262_gl_ram_ram_55_2 : DEL1BWP7T port map(I => gl_ram_ram_55(2), Z => FE_PHN262_gl_ram_ram_55_2);
  FE_PHC261_gl_ram_ram_54_1 : DEL1BWP7T port map(I => gl_ram_ram_54(1), Z => FE_PHN261_gl_ram_ram_54_1);
  FE_PHC260_gl_ram_ram_45_1 : DEL1BWP7T port map(I => gl_ram_ram_45(1), Z => FE_PHN260_gl_ram_ram_45_1);
  FE_PHC259_gl_ram_ram_95_2 : DEL1BWP7T port map(I => gl_ram_ram_95(2), Z => FE_PHN259_gl_ram_ram_95_2);
  FE_PHC258_gl_ram_ram_30_1 : DEL1BWP7T port map(I => gl_ram_ram_30(1), Z => FE_PHN258_gl_ram_ram_30_1);
  FE_PHC257_gl_ram_ram_98_0 : DEL1BWP7T port map(I => gl_ram_ram_98(0), Z => FE_PHN257_gl_ram_ram_98_0);
  FE_PHC256_gl_ram_ram_99_0 : DEL1BWP7T port map(I => gl_ram_ram_99(0), Z => FE_PHN256_gl_ram_ram_99_0);
  FE_PHC255_gl_ram_ram_70_0 : DEL1BWP7T port map(I => gl_ram_ram_70(0), Z => FE_PHN255_gl_ram_ram_70_0);
  FE_PHC254_gl_ram_ram_63_2 : DEL1BWP7T port map(I => gl_ram_ram_63(2), Z => FE_PHN254_gl_ram_ram_63_2);
  FE_PHC253_gl_ram_ram_61_0 : DEL1BWP7T port map(I => gl_ram_ram_61(0), Z => FE_PHN253_gl_ram_ram_61_0);
  FE_PHC252_gl_ram_ram_64_2 : DEL1BWP7T port map(I => gl_ram_ram_64(2), Z => FE_PHN252_gl_ram_ram_64_2);
  FE_PHC251_gl_ram_ram_28_0 : DEL1BWP7T port map(I => gl_ram_ram_28(0), Z => FE_PHN251_gl_ram_ram_28_0);
  FE_PHC250_gl_ram_ram_69_2 : DEL1BWP7T port map(I => gl_ram_ram_69(2), Z => FE_PHN250_gl_ram_ram_69_2);
  FE_PHC249_gl_ram_ram_55_0 : DEL1BWP7T port map(I => gl_ram_ram_55(0), Z => FE_PHN249_gl_ram_ram_55_0);
  FE_PHC248_gl_ram_ram_99_1 : DEL1BWP7T port map(I => gl_ram_ram_99(1), Z => FE_PHN248_gl_ram_ram_99_1);
  FE_PHC247_gl_ram_ram_58_2 : DEL1BWP7T port map(I => gl_ram_ram_58(2), Z => FE_PHN247_gl_ram_ram_58_2);
  FE_PHC246_gl_ram_ram_74_1 : DEL1BWP7T port map(I => gl_ram_ram_74(1), Z => FE_PHN246_gl_ram_ram_74_1);
  FE_PHC245_gl_ram_ram_20_0 : DEL1BWP7T port map(I => gl_ram_ram_20(0), Z => FE_PHN245_gl_ram_ram_20_0);
  FE_PHC244_gl_ram_ram_61_2 : DEL1BWP7T port map(I => gl_ram_ram_61(2), Z => FE_PHN244_gl_ram_ram_61_2);
  FE_PHC243_gl_ram_ram_4_1 : DEL1BWP7T port map(I => gl_ram_ram_4(1), Z => FE_PHN243_gl_ram_ram_4_1);
  FE_PHC242_gl_ram_ram_81_2 : DEL1BWP7T port map(I => gl_ram_ram_81(2), Z => FE_PHN242_gl_ram_ram_81_2);
  FE_PHC241_gl_ram_ram_90_2 : DEL1BWP7T port map(I => gl_ram_ram_90(2), Z => FE_PHN241_gl_ram_ram_90_2);
  FE_PHC240_gl_ram_ram_78_2 : DEL1BWP7T port map(I => gl_ram_ram_78(2), Z => FE_PHN240_gl_ram_ram_78_2);
  FE_PHC239_gl_ram_ram_34_2 : DEL1BWP7T port map(I => gl_ram_ram_34(2), Z => FE_PHN239_gl_ram_ram_34_2);
  FE_PHC238_gl_ram_ram_79_2 : DEL1BWP7T port map(I => gl_ram_ram_79(2), Z => FE_PHN238_gl_ram_ram_79_2);
  FE_PHC237_gl_ram_ram_29_2 : DEL1BWP7T port map(I => gl_ram_ram_29(2), Z => FE_PHN237_gl_ram_ram_29_2);
  FE_PHC236_gl_ram_ram_85_1 : DEL1BWP7T port map(I => gl_ram_ram_85(1), Z => FE_PHN236_gl_ram_ram_85_1);
  FE_PHC235_gl_ram_ram_89_2 : DEL1BWP7T port map(I => gl_ram_ram_89(2), Z => FE_PHN235_gl_ram_ram_89_2);
  FE_PHC234_gl_ram_ram_74_2 : DEL1BWP7T port map(I => gl_ram_ram_74(2), Z => FE_PHN234_gl_ram_ram_74_2);
  FE_PHC233_gl_ram_ram_94_0 : DEL1BWP7T port map(I => gl_ram_ram_94(0), Z => FE_PHN233_gl_ram_ram_94_0);
  FE_PHC232_gl_ram_ram_62_1 : DEL1BWP7T port map(I => gl_ram_ram_62(1), Z => FE_PHN232_gl_ram_ram_62_1);
  FE_PHC231_gl_ram_ram_47_1 : DEL1BWP7T port map(I => gl_ram_ram_47(1), Z => FE_PHN231_gl_ram_ram_47_1);
  FE_PHC230_gl_ram_ram_84_1 : DEL1BWP7T port map(I => gl_ram_ram_84(1), Z => FE_PHN230_gl_ram_ram_84_1);
  FE_PHC229_gl_ram_ram_69_1 : DEL1BWP7T port map(I => gl_ram_ram_69(1), Z => FE_PHN229_gl_ram_ram_69_1);
  FE_PHC228_gl_ram_ram_59_0 : DEL1BWP7T port map(I => gl_ram_ram_59(0), Z => FE_PHN228_gl_ram_ram_59_0);
  FE_PHC227_gl_ram_ram_49_1 : DEL1BWP7T port map(I => gl_ram_ram_49(1), Z => FE_PHN227_gl_ram_ram_49_1);
  FE_PHC226_gl_ram_ram_77_2 : DEL1BWP7T port map(I => gl_ram_ram_77(2), Z => FE_PHN226_gl_ram_ram_77_2);
  FE_PHC225_gl_ram_ram_44_2 : DEL1BWP7T port map(I => gl_ram_ram_44(2), Z => FE_PHN225_gl_ram_ram_44_2);
  FE_PHC224_gl_ram_ram_95_1 : DEL1BWP7T port map(I => gl_ram_ram_95(1), Z => FE_PHN224_gl_ram_ram_95_1);
  FE_PHC223_gl_ram_ram_26_1 : DEL1BWP7T port map(I => gl_ram_ram_26(1), Z => FE_PHN223_gl_ram_ram_26_1);
  FE_PHC222_gl_ram_ram_41_1 : DEL1BWP7T port map(I => gl_ram_ram_41(1), Z => FE_PHN222_gl_ram_ram_41_1);
  FE_PHC221_gl_ram_ram_64_0 : DEL1BWP7T port map(I => gl_ram_ram_64(0), Z => FE_PHN221_gl_ram_ram_64_0);
  FE_PHC220_gl_ram_ram_93_0 : DEL1BWP7T port map(I => gl_ram_ram_93(0), Z => FE_PHN220_gl_ram_ram_93_0);
  FE_PHC219_gl_ram_ram_81_1 : DEL1BWP7T port map(I => gl_ram_ram_81(1), Z => FE_PHN219_gl_ram_ram_81_1);
  FE_PHC218_gl_ram_ram_26_2 : DEL1BWP7T port map(I => gl_ram_ram_26(2), Z => FE_PHN218_gl_ram_ram_26_2);
  FE_PHC217_gl_ram_ram_32_2 : DEL1BWP7T port map(I => gl_ram_ram_32(2), Z => FE_PHN217_gl_ram_ram_32_2);
  FE_PHC216_gl_ram_ram_89_1 : DEL1BWP7T port map(I => gl_ram_ram_89(1), Z => FE_PHN216_gl_ram_ram_89_1);
  FE_PHC215_gl_ram_ram_69_0 : DEL1BWP7T port map(I => gl_ram_ram_69(0), Z => FE_PHN215_gl_ram_ram_69_0);
  FE_PHC214_gl_ram_ram_98_1 : DEL1BWP7T port map(I => gl_ram_ram_98(1), Z => FE_PHN214_gl_ram_ram_98_1);
  FE_PHC213_gl_ram_ram_49_0 : DEL1BWP7T port map(I => gl_ram_ram_49(0), Z => FE_PHN213_gl_ram_ram_49_0);
  FE_PHC212_gl_ram_ram_75_1 : DEL1BWP7T port map(I => gl_ram_ram_75(1), Z => FE_PHN212_gl_ram_ram_75_1);
  FE_PHC211_gl_ram_ram_57_0 : DEL1BWP7T port map(I => gl_ram_ram_57(0), Z => FE_PHN211_gl_ram_ram_57_0);
  FE_PHC210_gl_ram_ram_96_0 : DEL1BWP7T port map(I => gl_ram_ram_96(0), Z => FE_PHN210_gl_ram_ram_96_0);
  FE_PHC209_gl_ram_ram_80_2 : DEL1BWP7T port map(I => gl_ram_ram_80(2), Z => FE_PHN209_gl_ram_ram_80_2);
  FE_PHC208_gl_ram_ram_49_2 : DEL1BWP7T port map(I => gl_ram_ram_49(2), Z => FE_PHN208_gl_ram_ram_49_2);
  FE_PHC207_gl_ram_ram_62_2 : DEL1BWP7T port map(I => gl_ram_ram_62(2), Z => FE_PHN207_gl_ram_ram_62_2);
  FE_PHC206_gl_ram_ram_47_2 : DEL1BWP7T port map(I => gl_ram_ram_47(2), Z => FE_PHN206_gl_ram_ram_47_2);
  FE_PHC205_gl_ram_ram_14_1 : DEL1BWP7T port map(I => gl_ram_ram_14(1), Z => FE_PHN205_gl_ram_ram_14_1);
  FE_PHC204_gl_ram_ram_15_0 : DEL1BWP7T port map(I => gl_ram_ram_15(0), Z => FE_PHN204_gl_ram_ram_15_0);
  FE_PHC203_gl_ram_ram_2_1 : DEL1BWP7T port map(I => gl_ram_ram_2(1), Z => FE_PHN203_gl_ram_ram_2_1);
  FE_PHC202_gl_ram_ram_38_2 : DEL1BWP7T port map(I => gl_ram_ram_38(2), Z => FE_PHN202_gl_ram_ram_38_2);
  FE_PHC201_gl_ram_ram_30_0 : DEL1BWP7T port map(I => gl_ram_ram_30(0), Z => FE_PHN201_gl_ram_ram_30_0);
  FE_PHC200_gl_ram_ram_67_1 : DEL1BWP7T port map(I => gl_ram_ram_67(1), Z => FE_PHN200_gl_ram_ram_67_1);
  FE_PHC199_gl_ram_ram_77_1 : DEL1BWP7T port map(I => gl_ram_ram_77(1), Z => FE_PHN199_gl_ram_ram_77_1);
  FE_PHC198_gl_ram_ram_54_2 : DEL1BWP7T port map(I => gl_ram_ram_54(2), Z => FE_PHN198_gl_ram_ram_54_2);
  FE_PHC197_ml_il_y1_state_0 : DEL2BWP7T port map(I => FE_PHN197_ml_il_y1_state_0, Z => ml_il_y1_state(0));
  FE_PHC196_gl_ram_ram_72_2 : DEL1BWP7T port map(I => gl_ram_ram_72(2), Z => FE_PHN196_gl_ram_ram_72_2);
  FE_PHC195_gl_ram_ram_7_0 : DEL1BWP7T port map(I => gl_ram_ram_7(0), Z => FE_PHN195_gl_ram_ram_7_0);
  FE_PHC194_gl_ram_ram_1_1 : DEL1BWP7T port map(I => gl_ram_ram_1(1), Z => FE_PHN194_gl_ram_ram_1_1);
  FE_PHC193_gl_ram_ram_90_1 : DEL1BWP7T port map(I => gl_ram_ram_90(1), Z => FE_PHN193_gl_ram_ram_90_1);
  FE_PHC192_gl_ram_ram_16_0 : DEL1BWP7T port map(I => gl_ram_ram_16(0), Z => FE_PHN192_gl_ram_ram_16_0);
  FE_PHC191_gl_ram_ram_75_2 : DEL1BWP7T port map(I => gl_ram_ram_75(2), Z => FE_PHN191_gl_ram_ram_75_2);
  FE_PHC190_gl_ram_ram_93_1 : DEL1BWP7T port map(I => gl_ram_ram_93(1), Z => FE_PHN190_gl_ram_ram_93_1);
  FE_PHC189_gl_ram_ram_76_1 : DEL1BWP7T port map(I => gl_ram_ram_76(1), Z => FE_PHN189_gl_ram_ram_76_1);
  FE_PHC188_gl_ram_ram_83_2 : DEL1BWP7T port map(I => gl_ram_ram_83(2), Z => FE_PHN188_gl_ram_ram_83_2);
  FE_PHC187_gl_ram_ram_34_0 : DEL1BWP7T port map(I => gl_ram_ram_34(0), Z => FE_PHN187_gl_ram_ram_34_0);
  FE_PHC186_gl_ram_ram_30_2 : DEL1BWP7T port map(I => gl_ram_ram_30(2), Z => FE_PHN186_gl_ram_ram_30_2);
  FE_PHC185_gl_ram_ram_58_0 : DEL1BWP7T port map(I => gl_ram_ram_58(0), Z => FE_PHN185_gl_ram_ram_58_0);
  FE_PHC184_gl_ram_ram_21_1 : DEL1BWP7T port map(I => gl_ram_ram_21(1), Z => FE_PHN184_gl_ram_ram_21_1);
  FE_PHC183_gl_ram_ram_22_2 : DEL1BWP7T port map(I => gl_ram_ram_22(2), Z => FE_PHN183_gl_ram_ram_22_2);
  FE_PHC182_gl_ram_ram_25_2 : DEL1BWP7T port map(I => gl_ram_ram_25(2), Z => FE_PHN182_gl_ram_ram_25_2);
  FE_PHC181_gl_gr_lg_lh_n_17 : DEL1BWP7T port map(I => gl_gr_lg_lh_n_17, Z => FE_PHN181_gl_gr_lg_lh_n_17);
  FE_PHC180_gl_ram_ram_39_1 : DEL1BWP7T port map(I => gl_ram_ram_39(1), Z => FE_PHN180_gl_ram_ram_39_1);
  FE_PHC179_gl_ram_ram_51_0 : DEL1BWP7T port map(I => gl_ram_ram_51(0), Z => FE_PHN179_gl_ram_ram_51_0);
  FE_PHC178_gl_ram_ram_52_0 : DEL1BWP7T port map(I => gl_ram_ram_52(0), Z => FE_PHN178_gl_ram_ram_52_0);
  FE_PHC177_gl_ram_ram_13_2 : DEL1BWP7T port map(I => gl_ram_ram_13(2), Z => FE_PHN177_gl_ram_ram_13_2);
  FE_PHC176_gl_ram_ram_26_0 : DEL1BWP7T port map(I => gl_ram_ram_26(0), Z => FE_PHN176_gl_ram_ram_26_0);
  FE_PHC175_gl_ram_ram_15_1 : DEL1BWP7T port map(I => gl_ram_ram_15(1), Z => FE_PHN175_gl_ram_ram_15_1);
  FE_PHC174_gl_ram_ram_31_1 : DEL1BWP7T port map(I => gl_ram_ram_31(1), Z => FE_PHN174_gl_ram_ram_31_1);
  FE_PHC173_gl_ram_ram_7_1 : DEL1BWP7T port map(I => gl_ram_ram_7(1), Z => FE_PHN173_gl_ram_ram_7_1);
  FE_PHC172_gl_ram_ram_31_0 : DEL1BWP7T port map(I => gl_ram_ram_31(0), Z => FE_PHN172_gl_ram_ram_31_0);
  FE_PHC171_gl_ram_ram_3_1 : DEL1BWP7T port map(I => gl_ram_ram_3(1), Z => FE_PHN171_gl_ram_ram_3_1);
  FE_PHC170_ml_il_x1_state_0 : DEL1BWP7T port map(I => FE_PHN170_ml_il_x1_state_0, Z => ml_il_x1_state(0));
  FE_PHC169_gl_ram_ram_35_1 : DEL1BWP7T port map(I => gl_ram_ram_35(1), Z => FE_PHN169_gl_ram_ram_35_1);
  FE_PHC168_gl_ram_ram_91_0 : DEL1BWP7T port map(I => gl_ram_ram_91(0), Z => FE_PHN168_gl_ram_ram_91_0);
  FE_PHC167_gl_ram_ram_42_0 : DEL1BWP7T port map(I => gl_ram_ram_42(0), Z => FE_PHN167_gl_ram_ram_42_0);
  FE_PHC166_gl_ram_ram_10_2 : DEL1BWP7T port map(I => gl_ram_ram_10(2), Z => FE_PHN166_gl_ram_ram_10_2);
  FE_PHC165_gl_ram_ram_48_0 : DEL1BWP7T port map(I => gl_ram_ram_48(0), Z => FE_PHN165_gl_ram_ram_48_0);
  FE_PHC164_gl_ram_ram_91_2 : DEL1BWP7T port map(I => gl_ram_ram_91(2), Z => FE_PHN164_gl_ram_ram_91_2);
  FE_PHC163_gl_ram_ram_40_2 : DEL1BWP7T port map(I => gl_ram_ram_40(2), Z => FE_PHN163_gl_ram_ram_40_2);
  FE_PHC162_gl_ram_ram_74_0 : DEL1BWP7T port map(I => gl_ram_ram_74(0), Z => FE_PHN162_gl_ram_ram_74_0);
  FE_PHC161_gl_ram_ram_85_0 : DEL1BWP7T port map(I => gl_ram_ram_85(0), Z => FE_PHN161_gl_ram_ram_85_0);
  FE_PHC160_gl_ram_ram_10_1 : DEL1BWP7T port map(I => gl_ram_ram_10(1), Z => FE_PHN160_gl_ram_ram_10_1);
  FE_PHC159_gl_ram_ram_92_0 : DEL1BWP7T port map(I => gl_ram_ram_92(0), Z => FE_PHN159_gl_ram_ram_92_0);
  FE_PHC158_gl_ram_ram_19_2 : DEL1BWP7T port map(I => gl_ram_ram_19(2), Z => FE_PHN158_gl_ram_ram_19_2);
  FE_PHC157_gl_ram_ram_70_1 : DEL1BWP7T port map(I => gl_ram_ram_70(1), Z => FE_PHN157_gl_ram_ram_70_1);
  FE_PHC156_gl_ram_ram_94_2 : DEL1BWP7T port map(I => gl_ram_ram_94(2), Z => FE_PHN156_gl_ram_ram_94_2);
  FE_PHC155_gl_ram_ram_23_0 : DEL1BWP7T port map(I => gl_ram_ram_23(0), Z => FE_PHN155_gl_ram_ram_23_0);
  FE_PHC154_gl_ram_ram_84_0 : DEL1BWP7T port map(I => gl_ram_ram_84(0), Z => FE_PHN154_gl_ram_ram_84_0);
  FE_PHC153_gl_ram_ram_83_1 : DEL1BWP7T port map(I => gl_ram_ram_83(1), Z => FE_PHN153_gl_ram_ram_83_1);
  FE_PHC152_gl_ram_ram_79_0 : DEL1BWP7T port map(I => gl_ram_ram_79(0), Z => FE_PHN152_gl_ram_ram_79_0);
  FE_PHC151_gl_ram_ram_28_2 : DEL1BWP7T port map(I => gl_ram_ram_28(2), Z => FE_PHN151_gl_ram_ram_28_2);
  FE_PHC150_gl_ram_ram_81_0 : DEL1BWP7T port map(I => gl_ram_ram_81(0), Z => FE_PHN150_gl_ram_ram_81_0);
  FE_PHC149_gl_ram_ram_9_1 : DEL1BWP7T port map(I => gl_ram_ram_9(1), Z => FE_PHN149_gl_ram_ram_9_1);
  FE_PHC148_gl_ram_ram_56_0 : DEL1BWP7T port map(I => gl_ram_ram_56(0), Z => FE_PHN148_gl_ram_ram_56_0);
  FE_PHC147_gl_ram_ram_90_0 : DEL1BWP7T port map(I => gl_ram_ram_90(0), Z => FE_PHN147_gl_ram_ram_90_0);
  FE_PHC146_gl_ram_ram_38_0 : DEL1BWP7T port map(I => gl_ram_ram_38(0), Z => FE_PHN146_gl_ram_ram_38_0);
  FE_PHC145_gl_ram_ram_45_2 : DEL1BWP7T port map(I => gl_ram_ram_45(2), Z => FE_PHN145_gl_ram_ram_45_2);
  FE_PHC144_gl_ram_ram_65_1 : DEL1BWP7T port map(I => gl_ram_ram_65(1), Z => FE_PHN144_gl_ram_ram_65_1);
  FE_PHC143_gl_ram_ram_66_1 : DEL1BWP7T port map(I => gl_ram_ram_66(1), Z => FE_PHN143_gl_ram_ram_66_1);
  FE_PHC142_gl_ram_ram_93_2 : DEL1BWP7T port map(I => gl_ram_ram_93(2), Z => FE_PHN142_gl_ram_ram_93_2);
  FE_PHC141_gl_ram_ram_78_0 : DEL1BWP7T port map(I => gl_ram_ram_78(0), Z => FE_PHN141_gl_ram_ram_78_0);
  FE_PHC140_gl_ram_ram_12_0 : DEL1BWP7T port map(I => gl_ram_ram_12(0), Z => FE_PHN140_gl_ram_ram_12_0);
  FE_PHC139_gl_ram_ram_72_1 : DEL1BWP7T port map(I => gl_ram_ram_72(1), Z => FE_PHN139_gl_ram_ram_72_1);
  FE_PHC138_gl_ram_ram_46_0 : DEL1BWP7T port map(I => gl_ram_ram_46(0), Z => FE_PHN138_gl_ram_ram_46_0);
  FE_PHC137_gl_ram_ram_28_1 : DEL1BWP7T port map(I => gl_ram_ram_28(1), Z => FE_PHN137_gl_ram_ram_28_1);
  FE_PHC136_gl_ram_ram_18_1 : DEL1BWP7T port map(I => gl_ram_ram_18(1), Z => FE_PHN136_gl_ram_ram_18_1);
  FE_PHC135_gl_ram_ram_79_1 : DEL1BWP7T port map(I => gl_ram_ram_79(1), Z => FE_PHN135_gl_ram_ram_79_1);
  FE_PHC134_gl_ram_ram_57_2 : DEL1BWP7T port map(I => gl_ram_ram_57(2), Z => FE_PHN134_gl_ram_ram_57_2);
  FE_PHC133_gl_ram_ram_52_1 : DEL1BWP7T port map(I => gl_ram_ram_52(1), Z => FE_PHN133_gl_ram_ram_52_1);
  FE_PHC132_gl_ram_ram_80_1 : DEL1BWP7T port map(I => gl_ram_ram_80(1), Z => FE_PHN132_gl_ram_ram_80_1);
  FE_PHC131_gl_ram_ram_17_0 : DEL1BWP7T port map(I => gl_ram_ram_17(0), Z => FE_PHN131_gl_ram_ram_17_0);
  FE_PHC130_gl_ram_ram_71_0 : DEL1BWP7T port map(I => gl_ram_ram_71(0), Z => FE_PHN130_gl_ram_ram_71_0);
  FE_PHC129_gl_ram_ram_71_2 : DEL1BWP7T port map(I => gl_ram_ram_71(2), Z => FE_PHN129_gl_ram_ram_71_2);
  FE_PHC128_gl_ram_ram_68_1 : DEL1BWP7T port map(I => gl_ram_ram_68(1), Z => FE_PHN128_gl_ram_ram_68_1);
  FE_PHC127_gl_ram_ram_37_1 : DEL1BWP7T port map(I => gl_ram_ram_37(1), Z => FE_PHN127_gl_ram_ram_37_1);
  FE_PHC126_gl_ram_ram_13_1 : DEL1BWP7T port map(I => gl_ram_ram_13(1), Z => FE_PHN126_gl_ram_ram_13_1);
  FE_PHC125_gl_ram_ram_65_0 : DEL1BWP7T port map(I => gl_ram_ram_65(0), Z => FE_PHN125_gl_ram_ram_65_0);
  FE_PHC124_gl_ram_ram_62_0 : DEL1BWP7T port map(I => gl_ram_ram_62(0), Z => FE_PHN124_gl_ram_ram_62_0);
  FE_PHC123_ml_ms_count_debounce_11 : DEL1BWP7T port map(I => ml_ms_count_debounce(11), Z => FE_PHN123_ml_ms_count_debounce_11);
  FE_PHC122_gl_ram_ram_51_1 : DEL1BWP7T port map(I => gl_ram_ram_51(1), Z => FE_PHN122_gl_ram_ram_51_1);
  FE_PHC121_gl_ram_ram_50_0 : DEL1BWP7T port map(I => gl_ram_ram_50(0), Z => FE_PHN121_gl_ram_ram_50_0);
  FE_PHC120_gl_ram_ram_45_0 : DEL1BWP7T port map(I => gl_ram_ram_45(0), Z => FE_PHN120_gl_ram_ram_45_0);
  FE_PHC119_gl_ram_ram_29_0 : DEL1BWP7T port map(I => gl_ram_ram_29(0), Z => FE_PHN119_gl_ram_ram_29_0);
  FE_PHC118_gl_ram_ram_59_1 : DEL1BWP7T port map(I => gl_ram_ram_59(1), Z => FE_PHN118_gl_ram_ram_59_1);
  FE_PHC117_gl_ram_ram_53_2 : DEL1BWP7T port map(I => gl_ram_ram_53(2), Z => FE_PHN117_gl_ram_ram_53_2);
  FE_PHC116_gl_ram_ram_67_2 : DEL1BWP7T port map(I => gl_ram_ram_67(2), Z => FE_PHN116_gl_ram_ram_67_2);
  FE_PHC115_gl_ram_ram_95_0 : DEL1BWP7T port map(I => gl_ram_ram_95(0), Z => FE_PHN115_gl_ram_ram_95_0);
  FE_PHC114_gl_ram_ram_64_1 : DEL1BWP7T port map(I => gl_ram_ram_64(1), Z => FE_PHN114_gl_ram_ram_64_1);
  FE_PHC113_gl_ram_ram_99_2 : DEL1BWP7T port map(I => gl_ram_ram_99(2), Z => FE_PHN113_gl_ram_ram_99_2);
  FE_PHC112_gl_ram_ram_87_0 : DEL1BWP7T port map(I => gl_ram_ram_87(0), Z => FE_PHN112_gl_ram_ram_87_0);
  FE_PHC111_gl_ram_ram_44_1 : DEL1BWP7T port map(I => gl_ram_ram_44(1), Z => FE_PHN111_gl_ram_ram_44_1);
  FE_PHC110_gl_ram_ram_88_2 : DEL1BWP7T port map(I => gl_ram_ram_88(2), Z => FE_PHN110_gl_ram_ram_88_2);
  FE_PHC109_gl_ram_ram_85_2 : DEL1BWP7T port map(I => gl_ram_ram_85(2), Z => FE_PHN109_gl_ram_ram_85_2);
  FE_PHC108_gl_ram_ram_92_2 : DEL1BWP7T port map(I => gl_ram_ram_92(2), Z => FE_PHN108_gl_ram_ram_92_2);
  FE_PHC107_gl_ram_ram_72_0 : DEL1BWP7T port map(I => gl_ram_ram_72(0), Z => FE_PHN107_gl_ram_ram_72_0);
  FE_PHC106_gl_ram_ram_94_1 : DEL1BWP7T port map(I => gl_ram_ram_94(1), Z => FE_PHN106_gl_ram_ram_94_1);
  FE_PHC105_gl_ram_ram_21_2 : DEL1BWP7T port map(I => gl_ram_ram_21(2), Z => FE_PHN105_gl_ram_ram_21_2);
  FE_PHC104_gl_ram_ram_88_1 : DEL1BWP7T port map(I => gl_ram_ram_88(1), Z => FE_PHN104_gl_ram_ram_88_1);
  FE_PHC103_gl_ram_ram_68_2 : DEL1BWP7T port map(I => gl_ram_ram_68(2), Z => FE_PHN103_gl_ram_ram_68_2);
  FE_PHC102_gl_ram_ram_5_2 : DEL1BWP7T port map(I => gl_ram_ram_5(2), Z => FE_PHN102_gl_ram_ram_5_2);
  FE_PHC101_gl_ram_ram_92_1 : DEL1BWP7T port map(I => gl_ram_ram_92(1), Z => FE_PHN101_gl_ram_ram_92_1);
  FE_PHC100_gl_ram_ram_54_0 : DEL1BWP7T port map(I => gl_ram_ram_54(0), Z => FE_PHN100_gl_ram_ram_54_0);
  FE_PHC99_gl_ram_ram_97_2 : DEL1BWP7T port map(I => gl_ram_ram_97(2), Z => FE_PHN99_gl_ram_ram_97_2);
  FE_PHC98_gl_ram_ram_77_0 : DEL1BWP7T port map(I => gl_ram_ram_77(0), Z => FE_PHN98_gl_ram_ram_77_0);
  FE_PHC97_gl_ram_ram_16_1 : DEL1BWP7T port map(I => gl_ram_ram_16(1), Z => FE_PHN97_gl_ram_ram_16_1);
  FE_PHC96_gl_ram_ram_17_2 : DEL1BWP7T port map(I => gl_ram_ram_17(2), Z => FE_PHN96_gl_ram_ram_17_2);
  FE_PHC95_gl_ram_ram_7_2 : DEL1BWP7T port map(I => gl_ram_ram_7(2), Z => FE_PHN95_gl_ram_ram_7_2);
  FE_PHC94_gl_ram_ram_4_2 : DEL1BWP7T port map(I => gl_ram_ram_4(2), Z => FE_PHN94_gl_ram_ram_4_2);
  FE_PHC93_gl_gr_lg_lh_n_15 : DEL1BWP7T port map(I => gl_gr_lg_lh_n_15, Z => FE_PHN93_gl_gr_lg_lh_n_15);
  FE_PHC92_gl_ram_ram_84_2 : DEL1BWP7T port map(I => gl_ram_ram_84(2), Z => FE_PHN92_gl_ram_ram_84_2);
  FE_PHC91_ml_ms_cnt_n_0 : DEL1BWP7T port map(I => ml_ms_cnt_n_0, Z => FE_PHN91_ml_ms_cnt_n_0);
  FE_PHC90_ml_ms_data_sr_11bit_4 : DEL1BWP7T port map(I => FE_PHN90_ml_ms_data_sr_11bit_4, Z => ml_ms_data_sr_11bit(4));
  FE_PHC89_ml_ms_cntD_n_0 : DEL1BWP7T port map(I => ml_ms_cntD_n_0, Z => FE_PHN89_ml_ms_cntD_n_0);
  FE_PHC88_gl_vga_buf_Vint : DEL1BWP7T port map(I => FE_PHN88_gl_vga_buf_Vint, Z => gl_vga_buf_Vint);
  FE_PHC87_ml_il_color1_state_hs_0 : DEL0BWP7T port map(I => ml_il_color1_state_hs(0), Z => FE_PHN87_ml_il_color1_state_hs_0);
  FE_PHC86_ml_ms_sr11_data_out_0_79 : DEL1BWP7T port map(I => ml_ms_sr11_data_out_0_79, Z => FE_PHN86_ml_ms_sr11_data_out_0_79);
  FE_PHC85_ml_mouseX_2 : DEL1BWP7T port map(I => ml_mouseX(2), Z => FE_PHN85_ml_mouseX_2);
  FE_PHC84_ml_mouseX_1 : DEL1BWP7T port map(I => ml_mouseX(1), Z => FE_PHN84_ml_mouseX_1);
  FE_PHC83_clk15k_in : DEL1BWP7T port map(I => clk15k_in, Z => FE_PHN83_clk15k_in);
  FE_PHC82_ml_mouseY_2 : DEL1BWP7T port map(I => ml_mouseY(2), Z => FE_PHN82_ml_mouseY_2);
  FE_PHC81_gl_vga_buf_Bint : DEL1BWP7T port map(I => gl_vga_buf_Bint, Z => FE_PHN81_gl_vga_buf_Bint);
  FE_PHC80_ml_ms_sr11_data_out_5_84 : DEL1BWP7T port map(I => ml_ms_sr11_data_out_5_84, Z => FE_PHN80_ml_ms_sr11_data_out_5_84);
  FE_PHC79_ml_mouseY_1 : DEL1BWP7T port map(I => ml_mouseY(1), Z => FE_PHN79_ml_mouseY_1);
  FE_PHC78_ml_ms_sr11_data_out_1_80 : DEL1BWP7T port map(I => ml_ms_sr11_data_out_1_80, Z => FE_PHN78_ml_ms_sr11_data_out_1_80);
  FE_PHC77_ml_ms_n_26 : DEL1BWP7T port map(I => FE_PHN77_ml_ms_n_26, Z => ml_ms_n_26);
  FE_PHC76_ml_mouseX_0 : DEL1BWP7T port map(I => ml_mouseX(0), Z => FE_PHN76_ml_mouseX_0);
  FE_PHC75_ml_ms_n_20 : DEL1BWP7T port map(I => FE_PHN75_ml_ms_n_20, Z => ml_ms_n_20);
  FE_PHC74_ml_ms_n_19 : DEL1BWP7T port map(I => FE_PHN74_ml_ms_n_19, Z => ml_ms_n_19);
  FE_PHC73_ml_ms_n_25 : DEL1BWP7T port map(I => FE_PHN73_ml_ms_n_25, Z => ml_ms_n_25);
  FE_PHC72_ml_ms_data_sr_11bit_6 : DEL1BWP7T port map(I => FE_PHN72_ml_ms_data_sr_11bit_6, Z => ml_ms_data_sr_11bit(6));
  FE_PHC71_gl_vga_buf_Rint : DEL1BWP7T port map(I => gl_vga_buf_Rint, Z => FE_PHN71_gl_vga_buf_Rint);
  FE_PHC70_gl_vga_buf_Hint : DEL1BWP7T port map(I => gl_vga_buf_Hint, Z => FE_PHN70_gl_vga_buf_Hint);
  FE_PHC69_ml_ms_count_debounce_5 : DEL1BWP7T port map(I => ml_ms_count_debounce(5), Z => FE_PHN69_ml_ms_count_debounce_5);
  FE_PHC68_ml_ms_count_debounce_reset : DEL0BWP7T port map(I => ml_ms_count_debounce_reset, Z => FE_PHN68_ml_ms_count_debounce_reset);
  FE_PHC67_gl_vga_buf_Gint : DEL1BWP7T port map(I => gl_vga_buf_Gint, Z => FE_PHN67_gl_vga_buf_Gint);
  FE_PHC66_gl_vgd_vertical_9 : DEL1BWP7T port map(I => gl_vgd_vertical(9), Z => FE_PHN66_gl_vgd_vertical_9);
  FE_PHC65_ml_ms_count_debounce_4 : DEL1BWP7T port map(I => FE_PHN65_ml_ms_count_debounce_4, Z => ml_ms_count_debounce(4));
  FE_PHC64_ml_ms_count_debounce_3 : DEL1BWP7T port map(I => FE_PHN64_ml_ms_count_debounce_3, Z => ml_ms_count_debounce(3));
  FE_PHC63_ml_ms_count25M_7 : DEL0BWP7T port map(I => ml_ms_count25M(7), Z => FE_PHN63_ml_ms_count25M_7);
  FE_PHC62_ml_ms_count_debounce_8 : DEL1BWP7T port map(I => FE_PHN62_ml_ms_count_debounce_8, Z => ml_ms_count_debounce(8));
  FE_PHC61_ml_ms_count_debounce_9 : DEL1BWP7T port map(I => ml_ms_count_debounce(9), Z => FE_PHN61_ml_ms_count_debounce_9);
  FE_PHC60_ml_ms_cntD_count_0 : DEL1BWP7T port map(I => ml_ms_cntD_count(0), Z => FE_PHN60_ml_ms_cntD_count_0);
  FE_PHC59_ml_il_color1_n_1 : DEL0BWP7T port map(I => ml_il_color1_n_1, Z => FE_PHN59_ml_il_color1_n_1);
  FE_PHC58_ml_ms_cntD_count_2 : DEL1BWP7T port map(I => FE_PHN58_ml_ms_cntD_count_2, Z => ml_ms_cntD_count(2));
  FE_PHC57_gl_vgd_vertical_counter_8 : DEL1BWP7T port map(I => gl_vgd_vertical_counter(8), Z => FE_PHN57_gl_vgd_vertical_counter_8);
  FE_PHC56_ml_il_x1_state_1 : DEL1BWP7T port map(I => ml_il_x1_state(1), Z => FE_PHN56_ml_il_x1_state_1);
  FE_PHC55_ml_buttons_mouse_4 : DEL1BWP7T port map(I => ml_buttons_mouse(4), Z => FE_PHN55_ml_buttons_mouse_4);
  FE_PHC54_ml_il_y1_state_1 : DEL1BWP7T port map(I => FE_PHN54_ml_il_y1_state_1, Z => ml_il_y1_state(1));
  FE_PHC53_ml_ms_ed_reg1 : DEL1BWP7T port map(I => ml_ms_ed_reg1, Z => FE_PHN53_ml_ms_ed_reg1);
  FE_PHC52_gl_gr_lg_lv_l_edge_reg1 : DEL1BWP7T port map(I => gl_gr_lg_lv_l_edge_reg1, Z => FE_PHN52_gl_gr_lg_lv_l_edge_reg1);
  FE_PHC51_gl_gr_lg_lh_l_edge_reg1 : DEL1BWP7T port map(I => gl_gr_lg_lh_l_edge_reg1, Z => FE_PHN51_gl_gr_lg_lh_l_edge_reg1);
  FE_PHC50_gl_gr_lg_le_new_count_e_0 : DEL1BWP7T port map(I => FE_PHN50_gl_gr_lg_le_new_count_e_0, Z => gl_gr_lg_le_new_count_e(0));
  FE_PHC49_gl_gr_lg_le_new_count_e_1 : DEL1BWP7T port map(I => FE_PHN49_gl_gr_lg_le_new_count_e_1, Z => gl_gr_lg_le_new_count_e(1));
  FE_PHC48_gl_gr_lg_le_new_count_e_7 : DEL1BWP7T port map(I => gl_gr_lg_le_new_count_e(7), Z => FE_PHN48_gl_gr_lg_le_new_count_e_7);
  FE_PHC47_gl_gr_lg_le_new_count_e_2 : DEL1BWP7T port map(I => gl_gr_lg_le_new_count_e(2), Z => FE_PHN47_gl_gr_lg_le_new_count_e_2);
  FE_PHC46_gl_gr_lg_le_new_count_e_4 : DEL1BWP7T port map(I => gl_gr_lg_le_new_count_e(4), Z => FE_PHN46_gl_gr_lg_le_new_count_e_4);
  FE_PHC45_gl_gr_lg_le_new_count_e_9 : DEL1BWP7T port map(I => gl_gr_lg_le_new_count_e(9), Z => FE_PHN45_gl_gr_lg_le_new_count_e_9);
  FE_PHC44_gl_gr_lg_le_new_count_e_3 : DEL1BWP7T port map(I => gl_gr_lg_le_new_count_e(3), Z => FE_PHN44_gl_gr_lg_le_new_count_e_3);
  FE_PHC43_gl_gr_lg_le_new_count_e_8 : DEL1BWP7T port map(I => gl_gr_lg_le_new_count_e(8), Z => FE_PHN43_gl_gr_lg_le_new_count_e_8);
  FE_PHC42_gl_gr_lg_le_new_count_e_5 : DEL1BWP7T port map(I => gl_gr_lg_le_new_count_e(5), Z => FE_PHN42_gl_gr_lg_le_new_count_e_5);
  FE_PHC41_gl_gr_lg_le_new_count_e_6 : DEL1BWP7T port map(I => gl_gr_lg_le_new_count_e(6), Z => FE_PHN41_gl_gr_lg_le_new_count_e_6);
  FE_OFC40_gl_ram_n_16 : BUFFD1P5BWP7T port map(I => FE_OFN39_gl_ram_n_16, Z => FE_OFN40_gl_ram_n_16);
  FE_OFC39_gl_ram_n_16 : BUFFD1P5BWP7T port map(I => FE_OFN38_gl_ram_n_16, Z => FE_OFN39_gl_ram_n_16);
  FE_OFC38_gl_ram_n_16 : BUFFD1P5BWP7T port map(I => FE_OFN37_gl_ram_n_16, Z => FE_OFN38_gl_ram_n_16);
  FE_OFC37_gl_ram_n_16 : BUFFD2BWP7T port map(I => gl_ram_n_16, Z => FE_OFN37_gl_ram_n_16);
  FE_OFC36_clk15k_switch : BUFFD5BWP7T port map(I => FE_OFN36_clk15k_switch, Z => clk15k_switch);
  FE_OFC35_reset : DEL01BWP7T port map(I => reset, Z => FE_OFN35_reset);
  FE_OFC34_R : BUFFD5BWP7T port map(I => FE_OFN34_R, Z => R);
  FE_OFC33_B : BUFFD5BWP7T port map(I => FE_OFN33_B, Z => B);
  FE_OFC32_G : BUFFD5BWP7T port map(I => FE_OFN32_G, Z => G);
  FE_OFC31_H : BUFFD5BWP7T port map(I => FE_OFN31_H, Z => H);
  FE_OFC30_V : BUFFD5BWP7T port map(I => FE_OFN30_V, Z => V);
  FE_OFC29_gl_rom_n_20 : BUFFD1P5BWP7T port map(I => FE_OFN28_gl_rom_n_20, Z => FE_OFN29_gl_rom_n_20);
  FE_OFC28_gl_rom_n_20 : BUFFD1P5BWP7T port map(I => FE_OFN27_gl_rom_n_20, Z => FE_OFN28_gl_rom_n_20);
  FE_OFC27_gl_rom_n_20 : BUFFD1P5BWP7T port map(I => gl_rom_n_20, Z => FE_OFN27_gl_rom_n_20);
  FE_OFC26_gl_rom_n_19 : DEL01BWP7T port map(I => FE_OFN24_gl_rom_n_19, Z => FE_OFN26_gl_rom_n_19);
  FE_OFC25_gl_rom_n_19 : BUFFD1P5BWP7T port map(I => FE_OFN24_gl_rom_n_19, Z => FE_OFN25_gl_rom_n_19);
  FE_OFC24_gl_rom_n_19 : BUFFD2BWP7T port map(I => gl_rom_n_19, Z => FE_OFN24_gl_rom_n_19);
  FE_OFC23_gl_rom_n_21 : INVD1BWP7T port map(I => FE_OFN21_gl_rom_n_21, ZN => FE_OFN23_gl_rom_n_21);
  FE_OFC22_gl_rom_n_21 : CKND2BWP7T port map(I => FE_OFN21_gl_rom_n_21, ZN => FE_OFN22_gl_rom_n_21);
  FE_OFC21_gl_rom_n_21 : INVD1BWP7T port map(I => FE_OFN20_gl_rom_n_21, ZN => FE_OFN21_gl_rom_n_21);
  FE_OFC20_gl_rom_n_21 : BUFFD1P5BWP7T port map(I => FE_OFN19_gl_rom_n_21, Z => FE_OFN20_gl_rom_n_21);
  FE_OFC19_gl_rom_n_21 : BUFFD1P5BWP7T port map(I => gl_rom_n_21, Z => FE_OFN19_gl_rom_n_21);
  FE_OFC18_gl_rom_n_15 : CKND2BWP7T port map(I => FE_OFN16_gl_rom_n_15, ZN => FE_OFN18_gl_rom_n_15);
  FE_OFC17_gl_rom_n_15 : INVD1BWP7T port map(I => FE_OFN16_gl_rom_n_15, ZN => FE_OFN17_gl_rom_n_15);
  FE_OFC16_gl_rom_n_15 : INVD1BWP7T port map(I => FE_OFN15_gl_rom_n_15, ZN => FE_OFN16_gl_rom_n_15);
  FE_OFC15_gl_rom_n_15 : BUFFD2BWP7T port map(I => FE_OFN14_gl_rom_n_15, Z => FE_OFN15_gl_rom_n_15);
  FE_OFC14_gl_rom_n_15 : BUFFD1P5BWP7T port map(I => gl_rom_n_15, Z => FE_OFN14_gl_rom_n_15);
  FE_OFC13_gl_rom_n_22 : BUFFD2BWP7T port map(I => FE_OFN11_gl_rom_n_22, Z => FE_OFN13_gl_rom_n_22);
  FE_OFC12_gl_rom_n_22 : BUFFD1P5BWP7T port map(I => gl_rom_n_22, Z => FE_OFN12_gl_rom_n_22);
  FE_OFC11_gl_rom_n_22 : BUFFD1P5BWP7T port map(I => gl_rom_n_22, Z => FE_OFN11_gl_rom_n_22);
  FE_OFC10_gl_rom_n_17 : BUFFD2BWP7T port map(I => FE_OFN9_gl_rom_n_17, Z => FE_OFN10_gl_rom_n_17);
  FE_OFC9_gl_rom_n_17 : BUFFD2BWP7T port map(I => FE_OFN8_gl_rom_n_17, Z => FE_OFN9_gl_rom_n_17);
  FE_OFC8_gl_rom_n_17 : BUFFD2BWP7T port map(I => gl_rom_n_17, Z => FE_OFN8_gl_rom_n_17);
  FE_OFC7_gl_rom_n_18 : BUFFD1P5BWP7T port map(I => FE_OFN6_gl_rom_n_18, Z => FE_OFN7_gl_rom_n_18);
  FE_OFC6_gl_rom_n_18 : BUFFD1P5BWP7T port map(I => FE_OFN5_gl_rom_n_18, Z => FE_OFN6_gl_rom_n_18);
  FE_OFC5_gl_rom_n_18 : BUFFD2BWP7T port map(I => gl_rom_n_18, Z => FE_OFN5_gl_rom_n_18);
  FE_OFC4_gl_rom_n_16 : INVD1BWP7T port map(I => FE_OFN2_gl_rom_n_16, ZN => FE_OFN4_gl_rom_n_16);
  FE_OFC3_gl_rom_n_16 : CKND2BWP7T port map(I => FE_OFN2_gl_rom_n_16, ZN => FE_OFN3_gl_rom_n_16);
  FE_OFC2_gl_rom_n_16 : INVD1BWP7T port map(I => FE_OFN1_gl_rom_n_16, ZN => FE_OFN2_gl_rom_n_16);
  FE_OFC1_gl_rom_n_16 : BUFFD2BWP7T port map(I => FE_OFN0_gl_rom_n_16, Z => FE_OFN1_gl_rom_n_16);
  FE_OFC0_gl_rom_n_16 : BUFFD2BWP7T port map(I => gl_rom_n_16, Z => FE_OFN0_gl_rom_n_16);
  CTS_ccl_a_BUF_clk_G0_L2_5 : CKBD10BWP7T port map(I => CTS_24, Z => CTS_23);
  CTS_ccl_a_BUF_clk_G0_L2_4 : CKBD10BWP7T port map(I => CTS_24, Z => CTS_22);
  CTS_ccl_a_BUF_clk_G0_L2_3 : CKBD10BWP7T port map(I => CTS_24, Z => CTS_21);
  CTS_ccl_a_BUF_clk_G0_L2_2 : CKBD10BWP7T port map(I => CTS_24, Z => CTS_20);
  CTS_ccl_a_BUF_clk_G0_L2_1 : CKBD10BWP7T port map(I => CTS_24, Z => CTS_19);
  CTS_ccl_a_BUF_clk_G0_L1_1 : CKBD10BWP7T port map(I => clk, Z => CTS_24);
  FE_DBTC0_reset : INVD2BWP7T port map(I => FE_OFN35_reset, ZN => FE_DBTN0_reset);
  ml_il_x1_g901 : HA1D0BWP7T port map(A => ml_il_x1_input_register(3), B => ml_il_x1_n_27, CO => ml_il_x1_n_43, S => ml_il_x1_n_46);
  ml_il_x1_g902 : AO21D0BWP7T port map(A1 => ml_il_x1_n_28, A2 => ml_il_x1_input_register(3), B => ml_il_x1_n_44, Z => ml_il_x1_n_49);
  ml_il_x1_g903 : NR2D0BWP7T port map(A1 => ml_il_x1_n_28, A2 => ml_il_x1_input_register(3), ZN => ml_il_x1_n_44);
  ml_il_x1_g904 : OAI21D0BWP7T port map(A1 => ml_il_x1_n_26, A2 => ml_il_x1_n_21, B => ml_il_x1_n_22, ZN => ml_il_x1_n_28);
  ml_il_x1_g905 : MOAI22D0BWP7T port map(A1 => ml_il_x1_n_26, A2 => ml_il_x1_n_23, B1 => ml_il_x1_n_26, B2 => ml_il_x1_n_23, ZN => ml_il_x1_n_50);
  ml_il_x1_g906 : MOAI22D0BWP7T port map(A1 => ml_il_x1_n_25, A2 => ml_il_x1_n_20, B1 => ml_il_x1_input_register(2), B2 => ml_mouseX(2), ZN => ml_il_x1_n_27);
  ml_il_x1_g907 : CKXOR2D0BWP7T port map(A1 => ml_il_x1_n_23, A2 => ml_il_x1_n_25, Z => ml_il_x1_n_47);
  ml_il_x1_g908 : AOI21D0BWP7T port map(A1 => ml_il_x1_n_19, A2 => ml_il_x1_n_15, B => ml_il_x1_n_18, ZN => ml_il_x1_n_26);
  ml_il_x1_g909 : MOAI22D0BWP7T port map(A1 => ml_il_x1_n_24, A2 => ml_il_x1_n_16, B1 => ml_il_x1_n_24, B2 => ml_il_x1_n_16, ZN => ml_il_x1_n_48);
  ml_il_x1_g910 : MOAI22D0BWP7T port map(A1 => ml_il_x1_n_24, A2 => ml_il_x1_n_15, B1 => ml_il_x1_n_24, B2 => ml_il_x1_n_15, ZN => ml_il_x1_n_51);
  ml_il_x1_g911 : MAOI222D0BWP7T port map(A => ml_il_x1_input_register(1), B => ml_mouseX(1), C => ml_il_x1_n_17, ZN => ml_il_x1_n_25);
  ml_il_x1_g912 : IND2D0BWP7T port map(A1 => ml_il_x1_n_18, B1 => ml_il_x1_n_19, ZN => ml_il_x1_n_24);
  ml_il_x1_g913 : INR2D0BWP7T port map(A1 => ml_il_x1_n_22, B1 => ml_il_x1_n_21, ZN => ml_il_x1_n_23);
  ml_il_x1_g914 : NR2D0BWP7T port map(A1 => ml_il_x1_input_register(2), A2 => ml_mouseX(2), ZN => ml_il_x1_n_20);
  ml_il_x1_g915 : IND2D0BWP7T port map(A1 => ml_mouseX(2), B1 => ml_il_x1_input_register(2), ZN => ml_il_x1_n_22);
  ml_il_x1_g916 : INR2D0BWP7T port map(A1 => ml_mouseX(2), B1 => ml_il_x1_input_register(2), ZN => ml_il_x1_n_21);
  ml_il_x1_g917 : OAI21D0BWP7T port map(A1 => ml_il_x1_n_12, A2 => ml_mouseX(0), B => ml_il_x1_n_15, ZN => ml_il_x1_n_52);
  ml_il_x1_g918 : IND2D0BWP7T port map(A1 => ml_il_x1_input_register(1), B1 => ml_mouseX(1), ZN => ml_il_x1_n_19);
  ml_il_x1_g919 : INR2D0BWP7T port map(A1 => ml_il_x1_input_register(1), B1 => ml_mouseX(1), ZN => ml_il_x1_n_18);
  ml_il_x1_g920 : ND2D1BWP7T port map(A1 => ml_il_x1_n_13, A2 => FE_PHN395_ml_il_x1_n_9, ZN => ml_il_x1_input_register(2));
  ml_il_x1_g921 : ND2D1BWP7T port map(A1 => ml_il_x1_n_11, A2 => FE_PHN395_ml_il_x1_n_9, ZN => ml_il_x1_input_register(1));
  ml_il_x1_g922 : CKND1BWP7T port map(I => ml_il_x1_n_16, ZN => ml_il_x1_n_17);
  ml_il_x1_g923 : ND2D0BWP7T port map(A1 => ml_il_x1_input_register(0), A2 => ml_mouseX(0), ZN => ml_il_x1_n_16);
  ml_il_x1_g924 : ND2D0BWP7T port map(A1 => ml_il_x1_n_12, A2 => ml_mouseX(0), ZN => ml_il_x1_n_15);
  ml_il_x1_g925 : ND2D1BWP7T port map(A1 => ml_il_x1_n_14, A2 => FE_PHN395_ml_il_x1_n_9, ZN => ml_il_x1_input_register(3));
  ml_il_x1_g926 : AOI222D0BWP7T port map(A1 => ml_il_x1_n_10, A2 => ml_il_x1_n_46, B1 => ml_il_x1_n_7, B2 => ml_il_x1_n_49, C1 => ml_il_x1_n_5, C2 => sig_logic_x(3), ZN => ml_il_x1_n_14);
  ml_il_x1_g927 : AOI222D0BWP7T port map(A1 => ml_il_x1_n_10, A2 => ml_il_x1_n_47, B1 => ml_il_x1_n_7, B2 => ml_il_x1_n_50, C1 => ml_il_x1_n_5, C2 => sig_logic_x(2), ZN => ml_il_x1_n_13);
  ml_il_x1_g928 : INVD1BWP7T port map(I => ml_il_x1_n_12, ZN => ml_il_x1_input_register(0));
  ml_il_x1_g929 : AOI222D0BWP7T port map(A1 => ml_il_x1_n_10, A2 => ml_il_x1_n_48, B1 => ml_il_x1_n_7, B2 => ml_il_x1_n_51, C1 => ml_il_x1_n_5, C2 => sig_logic_x(1), ZN => ml_il_x1_n_11);
  ml_il_x1_g930 : AOI222D0BWP7T port map(A1 => ml_il_x1_n_10, A2 => ml_il_x1_n_52, B1 => ml_il_x1_n_7, B2 => ml_il_x1_n_52, C1 => ml_il_x1_n_5, C2 => sig_logic_x(0), ZN => ml_il_x1_n_12);
  ml_il_x1_g931 : NR3D0BWP7T port map(A1 => ml_il_x1_n_5, A2 => ml_buttons_mouse(0), A3 => ml_il_x1_n_8, ZN => ml_il_x1_n_10);
  ml_il_x1_g932 : IND3D1BWP7T port map(A1 => ml_buttons_mouse(0), B1 => ml_il_x1_n_8, B2 => ml_il_x1_state(0), ZN => ml_il_x1_n_9);
  ml_il_x1_g933 : IND2D0BWP7T port map(A1 => ml_il_x1_n_43, B1 => ml_il_x1_n_6, ZN => ml_il_x1_n_8);
  ml_il_x1_g934 : INR3D0BWP7T port map(A1 => ml_buttons_mouse(0), B1 => ml_il_x1_n_44, B2 => ml_il_x1_n_5, ZN => ml_il_x1_n_7);
  ml_il_x1_g935 : ND4D0BWP7T port map(A1 => ml_il_x1_n_47, A2 => ml_il_x1_n_48, A3 => ml_il_x1_n_52, A4 => ml_il_x1_n_46, ZN => ml_il_x1_n_6);
  ml_il_x1_state_reg_1 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => ml_il_x1_n_1, Q => ml_il_x1_state(1));
  ml_il_x1_g385 : INR4D0BWP7T port map(A1 => ml_handshake_mouse_out, B1 => FE_OFN35_reset, B2 => ml_il_x1_state(0), B3 => FE_PHN56_ml_il_x1_state_1, ZN => ml_il_x1_n_2);
  ml_il_x1_tempx_reg_0 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => ml_il_x1_input_register(0), Q => FE_PHN351_sig_logic_x_0);
  ml_il_x1_tempx_reg_1 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => ml_il_x1_input_register(1), Q => sig_logic_x(1));
  ml_il_x1_tempx_reg_2 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => ml_il_x1_input_register(2), Q => sig_logic_x(2));
  ml_il_x1_tempx_reg_3 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => ml_il_x1_input_register(3), Q => sig_logic_x(3));
  ml_il_x1_g390 : AO21D0BWP7T port map(A1 => ml_handshake_mouse_out, A2 => FE_PHN56_ml_il_x1_state_1, B => ml_il_x1_state(0), Z => ml_il_x1_n_1);
  ml_il_x1_state_reg_0 : DFD1BWP7T port map(CP => CTS_20, D => ml_il_x1_n_2, Q => FE_PHN170_ml_il_x1_state_0, QN => ml_il_x1_n_5);
  ml_il_y1_g901 : HA1D0BWP7T port map(A => ml_il_y1_input_register(3), B => ml_il_y1_n_27, CO => ml_il_y1_n_43, S => ml_il_y1_n_46);
  ml_il_y1_g902 : AO21D0BWP7T port map(A1 => ml_il_y1_n_28, A2 => ml_il_y1_input_register(3), B => ml_il_y1_n_44, Z => ml_il_y1_n_49);
  ml_il_y1_g903 : NR2D0BWP7T port map(A1 => ml_il_y1_n_28, A2 => ml_il_y1_input_register(3), ZN => ml_il_y1_n_44);
  ml_il_y1_g904 : OAI21D0BWP7T port map(A1 => ml_il_y1_n_26, A2 => ml_il_y1_n_21, B => ml_il_y1_n_22, ZN => ml_il_y1_n_28);
  ml_il_y1_g905 : MOAI22D0BWP7T port map(A1 => ml_il_y1_n_26, A2 => ml_il_y1_n_23, B1 => ml_il_y1_n_26, B2 => ml_il_y1_n_23, ZN => ml_il_y1_n_50);
  ml_il_y1_g906 : MOAI22D0BWP7T port map(A1 => ml_il_y1_n_25, A2 => ml_il_y1_n_20, B1 => ml_il_y1_input_register(2), B2 => ml_mouseY(2), ZN => ml_il_y1_n_27);
  ml_il_y1_g907 : CKXOR2D0BWP7T port map(A1 => ml_il_y1_n_23, A2 => ml_il_y1_n_25, Z => ml_il_y1_n_47);
  ml_il_y1_g908 : AOI21D0BWP7T port map(A1 => ml_il_y1_n_19, A2 => ml_il_y1_n_15, B => ml_il_y1_n_18, ZN => ml_il_y1_n_26);
  ml_il_y1_g909 : MOAI22D0BWP7T port map(A1 => ml_il_y1_n_24, A2 => ml_il_y1_n_16, B1 => ml_il_y1_n_24, B2 => ml_il_y1_n_16, ZN => ml_il_y1_n_48);
  ml_il_y1_g910 : MOAI22D0BWP7T port map(A1 => ml_il_y1_n_24, A2 => ml_il_y1_n_15, B1 => ml_il_y1_n_24, B2 => ml_il_y1_n_15, ZN => ml_il_y1_n_51);
  ml_il_y1_g911 : MAOI222D0BWP7T port map(A => ml_il_y1_input_register(1), B => ml_mouseY(1), C => ml_il_y1_n_17, ZN => ml_il_y1_n_25);
  ml_il_y1_g912 : IND2D0BWP7T port map(A1 => ml_il_y1_n_18, B1 => ml_il_y1_n_19, ZN => ml_il_y1_n_24);
  ml_il_y1_g913 : INR2D0BWP7T port map(A1 => ml_il_y1_n_22, B1 => ml_il_y1_n_21, ZN => ml_il_y1_n_23);
  ml_il_y1_g914 : NR2D0BWP7T port map(A1 => ml_il_y1_input_register(2), A2 => ml_mouseY(2), ZN => ml_il_y1_n_20);
  ml_il_y1_g915 : IND2D0BWP7T port map(A1 => ml_mouseY(2), B1 => ml_il_y1_input_register(2), ZN => ml_il_y1_n_22);
  ml_il_y1_g916 : INR2D0BWP7T port map(A1 => ml_mouseY(2), B1 => ml_il_y1_input_register(2), ZN => ml_il_y1_n_21);
  ml_il_y1_g917 : OAI21D0BWP7T port map(A1 => ml_il_y1_n_12, A2 => ml_mouseY(0), B => ml_il_y1_n_15, ZN => ml_il_y1_n_52);
  ml_il_y1_g918 : IND2D0BWP7T port map(A1 => ml_il_y1_input_register(1), B1 => ml_mouseY(1), ZN => ml_il_y1_n_19);
  ml_il_y1_g919 : INR2D0BWP7T port map(A1 => ml_il_y1_input_register(1), B1 => ml_mouseY(1), ZN => ml_il_y1_n_18);
  ml_il_y1_g920 : ND2D1BWP7T port map(A1 => ml_il_y1_n_13, A2 => FE_PHN384_ml_il_y1_n_9, ZN => ml_il_y1_input_register(2));
  ml_il_y1_g921 : ND2D1BWP7T port map(A1 => ml_il_y1_n_11, A2 => FE_PHN384_ml_il_y1_n_9, ZN => ml_il_y1_input_register(1));
  ml_il_y1_g922 : CKND1BWP7T port map(I => ml_il_y1_n_16, ZN => ml_il_y1_n_17);
  ml_il_y1_g923 : ND2D0BWP7T port map(A1 => ml_il_y1_input_register(0), A2 => ml_mouseY(0), ZN => ml_il_y1_n_16);
  ml_il_y1_g924 : ND2D0BWP7T port map(A1 => ml_il_y1_n_12, A2 => ml_mouseY(0), ZN => ml_il_y1_n_15);
  ml_il_y1_g925 : ND2D1BWP7T port map(A1 => ml_il_y1_n_14, A2 => FE_PHN384_ml_il_y1_n_9, ZN => ml_il_y1_input_register(3));
  ml_il_y1_g926 : AOI222D0BWP7T port map(A1 => ml_il_y1_n_10, A2 => ml_il_y1_n_46, B1 => ml_il_y1_n_7, B2 => ml_il_y1_n_49, C1 => ml_il_y1_n_5, C2 => sig_logic_y(3), ZN => ml_il_y1_n_14);
  ml_il_y1_g927 : AOI222D0BWP7T port map(A1 => ml_il_y1_n_10, A2 => ml_il_y1_n_47, B1 => ml_il_y1_n_7, B2 => ml_il_y1_n_50, C1 => ml_il_y1_n_5, C2 => sig_logic_y(2), ZN => ml_il_y1_n_13);
  ml_il_y1_g928 : INVD1BWP7T port map(I => ml_il_y1_n_12, ZN => ml_il_y1_input_register(0));
  ml_il_y1_g929 : AOI222D0BWP7T port map(A1 => ml_il_y1_n_10, A2 => ml_il_y1_n_48, B1 => ml_il_y1_n_7, B2 => ml_il_y1_n_51, C1 => ml_il_y1_n_5, C2 => sig_logic_y(1), ZN => ml_il_y1_n_11);
  ml_il_y1_g930 : AOI222D0BWP7T port map(A1 => ml_il_y1_n_10, A2 => ml_il_y1_n_52, B1 => ml_il_y1_n_7, B2 => ml_il_y1_n_52, C1 => ml_il_y1_n_5, C2 => sig_logic_y(0), ZN => ml_il_y1_n_12);
  ml_il_y1_g931 : NR3D0BWP7T port map(A1 => ml_il_y1_n_5, A2 => ml_buttons_mouse(1), A3 => ml_il_y1_n_8, ZN => ml_il_y1_n_10);
  ml_il_y1_g932 : IND3D1BWP7T port map(A1 => ml_buttons_mouse(1), B1 => ml_il_y1_n_8, B2 => ml_il_y1_state(0), ZN => ml_il_y1_n_9);
  ml_il_y1_g933 : IND2D0BWP7T port map(A1 => ml_il_y1_n_43, B1 => ml_il_y1_n_6, ZN => ml_il_y1_n_8);
  ml_il_y1_g934 : INR3D0BWP7T port map(A1 => ml_buttons_mouse(1), B1 => ml_il_y1_n_44, B2 => ml_il_y1_n_5, ZN => ml_il_y1_n_7);
  ml_il_y1_g935 : ND4D0BWP7T port map(A1 => ml_il_y1_n_47, A2 => ml_il_y1_n_48, A3 => ml_il_y1_n_52, A4 => ml_il_y1_n_46, ZN => ml_il_y1_n_6);
  ml_il_y1_state_reg_1 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_20, D => ml_il_y1_n_1, Q => FE_PHN54_ml_il_y1_state_1);
  ml_il_y1_g385 : INR4D0BWP7T port map(A1 => ml_handshake_mouse_out, B1 => FE_OFN35_reset, B2 => ml_il_y1_state(0), B3 => ml_il_y1_state(1), ZN => ml_il_y1_n_2);
  ml_il_y1_tempy_reg_0 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_20, D => ml_il_y1_input_register(0), Q => FE_PHN349_sig_logic_y_0);
  ml_il_y1_tempy_reg_1 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_20, D => ml_il_y1_input_register(1), Q => sig_logic_y(1));
  ml_il_y1_tempy_reg_2 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_20, D => ml_il_y1_input_register(2), Q => sig_logic_y(2));
  ml_il_y1_tempy_reg_3 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_20, D => ml_il_y1_input_register(3), Q => sig_logic_y(3));
  ml_il_y1_g390 : AO21D0BWP7T port map(A1 => ml_handshake_mouse_out, A2 => ml_il_y1_state(1), B => ml_il_y1_state(0), Z => ml_il_y1_n_1);
  ml_il_y1_state_reg_0 : DFD1BWP7T port map(CP => CTS_20, D => ml_il_y1_n_2, Q => FE_PHN197_ml_il_y1_state_0, QN => ml_il_y1_n_5);
  gl_gr_lg_x_grid_asked_reg_0 : LNQD1BWP7T port map(D => gl_n_62, EN => gl_n_66, Q => gl_sig_x(0));
  gl_gr_lg_x_grid_asked_reg_3 : LNQD1BWP7T port map(D => gl_n_59, EN => gl_n_66, Q => gl_sig_x(3));
  gl_gr_lg_y_grid_asked_reg_3 : LNQD1BWP7T port map(D => gl_n_58, EN => gl_n_66, Q => gl_sig_y(3));
  gl_gr_lg_y_grid_asked_reg_0 : LNQD1BWP7T port map(D => gl_n_60, EN => gl_n_66, Q => gl_sig_y(0));
  gl_gr_lg_y_grid_asked_reg_2 : LNQD1BWP7T port map(D => gl_n_57, EN => gl_n_66, Q => gl_sig_y(2));
  gl_gr_lg_x_grid_asked_reg_1 : LNQD1BWP7T port map(D => gl_n_56, EN => gl_n_66, Q => gl_sig_x(1));
  gl_gr_lg_x_grid_asked_reg_2 : LNQD1BWP7T port map(D => gl_n_61, EN => gl_n_66, Q => gl_sig_x(2));
  gl_gr_lg_y_grid_asked_reg_1 : LNQD1BWP7T port map(D => gl_n_55, EN => gl_n_66, Q => gl_sig_y(1));
  gl_g1441 : AOI21D0BWP7T port map(A1 => gl_n_65, A2 => gl_sig_rom(0), B => gl_n_64, ZN => gl_n_66);
  gl_g1442 : AOI21D0BWP7T port map(A1 => gl_n_63, A2 => gl_gr_lg_n_113, B => gl_sig_rom(1), ZN => gl_n_65);
  gl_g1443 : ND2D0BWP7T port map(A1 => gl_gr_lg_n_104, A2 => gl_n_53, ZN => gl_n_63);
  gl_g1444 : NR2D0BWP7T port map(A1 => gl_n_54, A2 => gl_gr_lg_local_x(0), ZN => gl_n_62);
  gl_g1445 : AOI21D0BWP7T port map(A1 => gl_n_45, A2 => gl_n_42, B => gl_n_54, ZN => gl_n_61);
  gl_g1446 : NR2D0BWP7T port map(A1 => gl_n_54, A2 => gl_gr_lg_local_y(0), ZN => gl_n_60);
  gl_g1447 : NR2D0BWP7T port map(A1 => gl_gr_lg_n_104, A2 => gl_gr_lg_n_113, ZN => gl_n_64);
  gl_g1448 : AN3D0BWP7T port map(A1 => gl_gr_lg_n_105, A2 => gl_n_45, A3 => gl_gr_lg_local_x(3), Z => gl_n_59);
  gl_g1449 : AN3D0BWP7T port map(A1 => gl_gr_lg_n_105, A2 => gl_n_46, A3 => gl_gr_lg_local_y(3), Z => gl_n_58);
  gl_g1450 : NR2D0BWP7T port map(A1 => gl_n_54, A2 => gl_n_47, ZN => gl_n_57);
  gl_g1451 : AOI21D0BWP7T port map(A1 => gl_n_35, A2 => gl_n_34, B => gl_n_54, ZN => gl_n_56);
  gl_g1452 : AOI21D0BWP7T port map(A1 => gl_n_33, A2 => gl_n_36, B => gl_n_54, ZN => gl_n_55);
  gl_g1454 : INVD1BWP7T port map(I => gl_n_54, ZN => gl_gr_lg_n_105);
  gl_g1455 : NR4D0BWP7T port map(A1 => gl_n_51, A2 => gl_n_40, A3 => gl_n_39, A4 => gl_n_43, ZN => gl_gr_lg_n_104);
  gl_g1456 : OAI211D1BWP7T port map(A1 => gl_gr_lg_local_y(3), A2 => gl_n_46, B => gl_n_52, C => gl_n_48, ZN => gl_n_54);
  gl_g1457 : NR4D0BWP7T port map(A1 => gl_n_49, A2 => gl_n_36, A3 => gl_gr_lg_local_y(2), A4 => gl_gr_lg_local_y(3), ZN => gl_gr_lg_n_113);
  gl_g1458 : CKND1BWP7T port map(I => gl_n_53, ZN => gl_n_52);
  gl_g1459 : NR2D1BWP7T port map(A1 => gl_n_45, A2 => gl_gr_lg_local_x(3), ZN => gl_n_53);
  gl_g1460 : ND4D0BWP7T port map(A1 => gl_n_50, A2 => gl_n_41, A3 => gl_n_38, A4 => gl_n_37, ZN => gl_n_51);
  gl_g1461 : AOI211XD0BWP7T port map(A1 => gl_n_29, A2 => sig_logic_x(3), B => gl_n_44, C => gl_n_32, ZN => gl_n_50);
  gl_g1462 : AN4D0BWP7T port map(A1 => gl_n_30, A2 => gl_gr_lg_local_x(2), A3 => gl_gr_lg_local_x(1), A4 => gl_gr_lg_local_x(3), Z => gl_n_49);
  gl_g1463 : AO21D0BWP7T port map(A1 => gl_n_34, A2 => gl_n_31, B => gl_n_29, Z => gl_n_48);
  gl_g1464 : XNR2D1BWP7T port map(A1 => gl_n_33, A2 => gl_gr_lg_local_y(2), ZN => gl_n_47);
  gl_g1465 : CKXOR2D1BWP7T port map(A1 => sig_logic_y(3), A2 => gl_gr_lg_local_y(3), Z => gl_n_44);
  gl_g1466 : MOAI22D0BWP7T port map(A1 => gl_n_31, A2 => sig_logic_x(2), B1 => gl_n_31, B2 => sig_logic_x(2), ZN => gl_n_43);
  gl_g1467 : ND2D0BWP7T port map(A1 => gl_n_35, A2 => gl_gr_lg_local_x(2), ZN => gl_n_42);
  gl_g1468 : CKAN2D1BWP7T port map(A1 => gl_n_33, A2 => gl_gr_lg_local_y(2), Z => gl_n_46);
  gl_g1469 : OR2D1BWP7T port map(A1 => gl_n_35, A2 => gl_gr_lg_local_x(2), Z => gl_n_45);
  gl_g1470 : XNR2D1BWP7T port map(A1 => sig_logic_y(2), A2 => gl_gr_lg_local_y(2), ZN => gl_n_41);
  gl_g1471 : CKXOR2D0BWP7T port map(A1 => gl_gr_lg_local_x(1), A2 => sig_logic_x(1), Z => gl_n_40);
  gl_g1472 : MOAI22D0BWP7T port map(A1 => gl_n_30, A2 => sig_logic_x(0), B1 => gl_n_30, B2 => sig_logic_x(0), ZN => gl_n_39);
  gl_g1473 : XNR2D1BWP7T port map(A1 => sig_logic_y(0), A2 => gl_gr_lg_local_y(0), ZN => gl_n_38);
  gl_g1474 : XNR2D1BWP7T port map(A1 => sig_logic_y(1), A2 => gl_gr_lg_local_y(1), ZN => gl_n_37);
  gl_g1475 : ND2D1BWP7T port map(A1 => gl_gr_lg_local_y(0), A2 => gl_gr_lg_local_y(1), ZN => gl_n_36);
  gl_g1476 : IND2D1BWP7T port map(A1 => gl_gr_lg_local_x(1), B1 => gl_n_30, ZN => gl_n_35);
  gl_g1477 : NR2D0BWP7T port map(A1 => gl_n_29, A2 => sig_logic_x(3), ZN => gl_n_32);
  gl_g1478 : CKND2D1BWP7T port map(A1 => gl_gr_lg_local_x(1), A2 => gl_gr_lg_local_x(0), ZN => gl_n_34);
  gl_g1479 : OR2D1BWP7T port map(A1 => gl_gr_lg_local_y(0), A2 => gl_gr_lg_local_y(1), Z => gl_n_33);
  gl_g1480 : INVD1BWP7T port map(I => gl_gr_lg_local_x(2), ZN => gl_n_31);
  gl_g1481 : INVD1BWP7T port map(I => gl_gr_lg_local_x(0), ZN => gl_n_30);
  gl_g1482 : INVD0BWP7T port map(I => gl_gr_lg_local_x(3), ZN => gl_n_29);
  gl_g1242 : ND4D0BWP7T port map(A1 => gl_n_28, A2 => gl_n_27, A3 => gl_n_11, A4 => gl_n_12, ZN => gl_sig_green);
  gl_g1243 : AOI222D0BWP7T port map(A1 => gl_n_25, A2 => gl_n_87, B1 => gl_n_21, B2 => gl_n_23, C1 => gl_n_26, C2 => gl_n_84, ZN => gl_n_28);
  gl_g1244 : MAOI22D0BWP7T port map(A1 => gl_n_4, A2 => sig_output_color(1), B1 => gl_n_16, B2 => gl_n_24, ZN => gl_n_27);
  gl_g1245 : AOI21D0BWP7T port map(A1 => gl_n_7, A2 => gl_n_2, B => gl_n_24, ZN => gl_n_26);
  gl_g1246 : AO32D1BWP7T port map(A1 => gl_n_22, A2 => gl_n_103, A3 => gl_gr_lg_local_x(3), B1 => gl_n_20, B2 => gl_n_23, Z => gl_n_25);
  gl_g1247 : IND3D1BWP7T port map(A1 => gl_n_87, B1 => gl_gr_lg_local_x(3), B2 => gl_n_23, ZN => gl_n_24);
  gl_g1248 : NR4D0BWP7T port map(A1 => gl_n_103, A2 => gl_n_102, A3 => gl_n_88, A4 => gl_n_126, ZN => gl_n_23);
  gl_g1249 : IINR4D0BWP7T port map(A1 => gl_n_102, A2 => gl_n_88, B1 => gl_n_19, B2 => gl_n_126, ZN => gl_n_22);
  gl_g1250 : OAI32D1BWP7T port map(A1 => gl_n_86, A2 => gl_n_0, A3 => gl_n_17, B1 => gl_n_87, B2 => gl_n_19, ZN => gl_n_21);
  gl_g1251 : MOAI22D0BWP7T port map(A1 => gl_n_16, A2 => gl_n_84, B1 => gl_n_3, B2 => gl_gr_lg_local_x(3), ZN => gl_n_20);
  gl_g1252 : ND2D1BWP7T port map(A1 => gl_n_11, A2 => gl_n_14, ZN => gl_sig_blue);
  gl_g1253 : ND2D1BWP7T port map(A1 => gl_n_11, A2 => gl_n_15, ZN => gl_sig_red);
  gl_g1254 : OAI21D0BWP7T port map(A1 => gl_n_8, A2 => gl_gr_lg_local_x(2), B => gl_n_87, ZN => gl_n_17);
  gl_g1255 : ND2D1BWP7T port map(A1 => gl_n_13, A2 => gl_gr_lg_local_x(2), ZN => gl_n_19);
  gl_g1257 : AOI22D0BWP7T port map(A1 => gl_n_9, A2 => gl_sig_ram(0), B1 => gl_n_4, B2 => sig_output_color(0), ZN => gl_n_15);
  gl_g1258 : AOI22D0BWP7T port map(A1 => gl_n_9, A2 => gl_sig_ram(2), B1 => gl_n_4, B2 => sig_output_color(2), ZN => gl_n_14);
  gl_g1259 : MAOI22D0BWP7T port map(A1 => gl_n_86, A2 => gl_gr_lg_local_x(2), B1 => gl_n_10, B2 => gl_n_2, ZN => gl_n_16);
  gl_g1260 : NR2D1BWP7T port map(A1 => gl_n_7, A2 => gl_n_3, ZN => gl_n_13);
  gl_g1261 : CKND2D0BWP7T port map(A1 => gl_n_9, A2 => gl_sig_ram(1), ZN => gl_n_12);
  gl_g1262 : INR2XD0BWP7T port map(A1 => gl_n_5, B1 => gl_gr_lg_local_x(1), ZN => gl_n_10);
  gl_g1263 : ND2D1BWP7T port map(A1 => gl_n_4, A2 => gl_sig_rom(0), ZN => gl_n_11);
  gl_g1264 : INVD1BWP7T port map(I => gl_n_7, ZN => gl_n_8);
  gl_g1266 : OA21D0BWP7T port map(A1 => gl_sig_rom(0), A2 => gl_n_1, B => gl_gr_lg_n_105, Z => gl_n_9);
  gl_g1267 : IND2D1BWP7T port map(A1 => gl_n_5, B1 => gl_gr_lg_local_x(1), ZN => gl_n_7);
  gl_g1268 : NR2XD0BWP7T port map(A1 => gl_n_85, A2 => gl_gr_lg_local_x(0), ZN => gl_n_5);
  gl_g1269 : AN2D1BWP7T port map(A1 => gl_sig_rom(1), A2 => gl_gr_lg_n_104, Z => gl_n_4);
  gl_g1270 : ND2D1BWP7T port map(A1 => gl_n_84, A2 => gl_n_86, ZN => gl_n_3);
  gl_g1271 : NR2XD0BWP7T port map(A1 => gl_n_86, A2 => gl_gr_lg_local_x(2), ZN => gl_n_2);
  gl_g1272 : INVD1BWP7T port map(I => gl_gr_lg_n_104, ZN => gl_n_1);
  gl_g1273 : INVD0BWP7T port map(I => gl_n_84, ZN => gl_n_0);
  gl_g2 : OAI21D0BWP7T port map(A1 => gl_n_125, A2 => gl_n_1, B => gl_gr_lg_n_113, ZN => gl_n_126);
  gl_g3 : INR2D1BWP7T port map(A1 => gl_sig_rom(0), B1 => gl_n_53, ZN => gl_n_125);
  gl_rom_rom_colour_out_reg_0 : LHQD1BWP7T port map(D => gl_rom_n_1500, E => CTS_19, Q => gl_sig_rom(0));
  gl_rom_rom_colour_out_reg_1 : LHQD1BWP7T port map(D => gl_rom_n_1499, E => CTS_19, Q => gl_sig_rom(1));
  gl_rom_g34917 : MOAI22D0BWP7T port map(A1 => gl_rom_n_1496, A2 => gl_sig_e(9), B1 => gl_rom_n_1498, B2 => gl_sig_e(9), ZN => gl_rom_n_1500);
  gl_rom_g34918 : MOAI22D0BWP7T port map(A1 => gl_rom_n_1497, A2 => gl_sig_e(9), B1 => gl_rom_n_1495, B2 => gl_sig_e(9), ZN => gl_rom_n_1499);
  gl_rom_g34919 : ND4D0BWP7T port map(A1 => gl_rom_n_1488, A2 => gl_rom_n_1480, A3 => gl_rom_n_1481, A4 => gl_rom_n_1490, ZN => gl_rom_n_1498);
  gl_rom_g34920 : AN4D0BWP7T port map(A1 => gl_rom_n_1484, A2 => gl_rom_n_1483, A3 => gl_rom_n_1482, A4 => gl_rom_n_1493, Z => gl_rom_n_1497);
  gl_rom_g34921 : AN4D0BWP7T port map(A1 => gl_rom_n_1485, A2 => gl_rom_n_1487, A3 => gl_rom_n_1494, A4 => gl_rom_n_1492, Z => gl_rom_n_1496);
  gl_rom_g34922 : ND4D0BWP7T port map(A1 => gl_rom_n_1486, A2 => gl_rom_n_1479, A3 => gl_rom_n_1489, A4 => gl_rom_n_1491, ZN => gl_rom_n_1495);
  gl_rom_g34923 : AOI22D0BWP7T port map(A1 => gl_rom_n_1475, A2 => gl_rom_n_33, B1 => gl_rom_n_1463, B2 => gl_rom_n_36, ZN => gl_rom_n_1494);
  gl_rom_g34924 : AOI22D0BWP7T port map(A1 => gl_rom_n_1472, A2 => gl_rom_n_37, B1 => gl_rom_n_1456, B2 => gl_rom_n_31, ZN => gl_rom_n_1493);
  gl_rom_g34925 : AOI22D0BWP7T port map(A1 => gl_rom_n_1460, A2 => gl_rom_n_37, B1 => gl_rom_n_1447, B2 => gl_rom_n_31, ZN => gl_rom_n_1492);
  gl_rom_g34926 : AOI22D0BWP7T port map(A1 => gl_rom_n_1477, A2 => gl_rom_n_37, B1 => gl_rom_n_1462, B2 => gl_rom_n_31, ZN => gl_rom_n_1491);
  gl_rom_g34927 : AOI22D0BWP7T port map(A1 => gl_rom_n_1458, A2 => gl_rom_n_37, B1 => gl_rom_n_1454, B2 => gl_rom_n_31, ZN => gl_rom_n_1490);
  gl_rom_g34928 : AOI22D0BWP7T port map(A1 => gl_rom_n_1474, A2 => gl_rom_n_32, B1 => gl_rom_n_1476, B2 => gl_rom_n_35, ZN => gl_rom_n_1489);
  gl_rom_g34929 : AOI22D0BWP7T port map(A1 => gl_rom_n_1452, A2 => gl_rom_n_32, B1 => gl_rom_n_1473, B2 => gl_rom_n_35, ZN => gl_rom_n_1488);
  gl_rom_g34930 : AOI22D0BWP7T port map(A1 => gl_rom_n_1470, A2 => gl_rom_n_38, B1 => gl_rom_n_1455, B2 => gl_rom_n_34, ZN => gl_rom_n_1487);
  gl_rom_g34931 : AOI22D0BWP7T port map(A1 => gl_rom_n_1449, A2 => gl_rom_n_33, B1 => gl_rom_n_1478, B2 => gl_rom_n_36, ZN => gl_rom_n_1486);
  gl_rom_g34932 : AOI22D0BWP7T port map(A1 => gl_rom_n_1465, A2 => gl_rom_n_32, B1 => gl_rom_n_1467, B2 => gl_rom_n_35, ZN => gl_rom_n_1485);
  gl_rom_g34933 : AOI22D0BWP7T port map(A1 => gl_rom_n_1466, A2 => gl_rom_n_33, B1 => gl_rom_n_1453, B2 => gl_rom_n_36, ZN => gl_rom_n_1484);
  gl_rom_g34934 : AOI22D0BWP7T port map(A1 => gl_rom_n_1464, A2 => gl_rom_n_32, B1 => gl_rom_n_1451, B2 => gl_rom_n_35, ZN => gl_rom_n_1483);
  gl_rom_g34935 : AOI22D0BWP7T port map(A1 => gl_rom_n_1468, A2 => gl_rom_n_38, B1 => gl_rom_n_1469, B2 => gl_rom_n_34, ZN => gl_rom_n_1482);
  gl_rom_g34936 : AOI22D0BWP7T port map(A1 => gl_rom_n_1471, A2 => gl_rom_n_33, B1 => gl_rom_n_1448, B2 => gl_rom_n_36, ZN => gl_rom_n_1481);
  gl_rom_g34937 : AOI22D0BWP7T port map(A1 => gl_rom_n_1457, A2 => gl_rom_n_38, B1 => gl_rom_n_1450, B2 => gl_rom_n_34, ZN => gl_rom_n_1480);
  gl_rom_g34938 : AOI22D0BWP7T port map(A1 => gl_rom_n_1459, A2 => gl_rom_n_38, B1 => gl_rom_n_1461, B2 => gl_rom_n_34, ZN => gl_rom_n_1479);
  gl_rom_g34939 : ND4D0BWP7T port map(A1 => gl_rom_n_1342, A2 => gl_rom_n_1424, A3 => gl_rom_n_1337, A4 => gl_rom_n_1340, ZN => gl_rom_n_1478);
  gl_rom_g34940 : ND4D0BWP7T port map(A1 => gl_rom_n_1407, A2 => gl_rom_n_1409, A3 => gl_rom_n_1445, A4 => gl_rom_n_1404, ZN => gl_rom_n_1477);
  gl_rom_g34941 : ND4D0BWP7T port map(A1 => gl_rom_n_1443, A2 => gl_rom_n_1398, A3 => gl_rom_n_1400, A4 => gl_rom_n_1403, ZN => gl_rom_n_1476);
  gl_rom_g34942 : ND4D0BWP7T port map(A1 => gl_rom_n_1401, A2 => gl_rom_n_1442, A3 => gl_rom_n_1396, A4 => gl_rom_n_1392, ZN => gl_rom_n_1475);
  gl_rom_g34943 : ND4D0BWP7T port map(A1 => gl_rom_n_1397, A2 => gl_rom_n_1394, A3 => gl_rom_n_1440, A4 => gl_rom_n_1391, ZN => gl_rom_n_1474);
  gl_rom_g34944 : ND4D0BWP7T port map(A1 => gl_rom_n_1435, A2 => gl_rom_n_1386, A3 => gl_rom_n_1381, A4 => gl_rom_n_1366, ZN => gl_rom_n_1473);
  gl_rom_g34945 : ND4D0BWP7T port map(A1 => gl_rom_n_1385, A2 => gl_rom_n_1437, A3 => gl_rom_n_1379, A4 => gl_rom_n_1383, ZN => gl_rom_n_1472);
  gl_rom_g34946 : ND4D0BWP7T port map(A1 => gl_rom_n_1350, A2 => gl_rom_n_1371, A3 => gl_rom_n_1427, A4 => gl_rom_n_1341, ZN => gl_rom_n_1471);
  gl_rom_g34947 : ND4D0BWP7T port map(A1 => gl_rom_n_1376, A2 => gl_rom_n_1434, A3 => gl_rom_n_1377, A4 => gl_rom_n_1368, ZN => gl_rom_n_1470);
  gl_rom_g34948 : ND4D0BWP7T port map(A1 => gl_rom_n_1378, A2 => gl_rom_n_1436, A3 => gl_rom_n_1374, A4 => gl_rom_n_1375, ZN => gl_rom_n_1469);
  gl_rom_g34949 : ND4D0BWP7T port map(A1 => gl_rom_n_1433, A2 => gl_rom_n_1369, A3 => gl_rom_n_1372, A4 => gl_rom_n_1370, ZN => gl_rom_n_1468);
  gl_rom_g34950 : ND4D0BWP7T port map(A1 => gl_rom_n_1365, A2 => gl_rom_n_1363, A3 => gl_rom_n_1357, A4 => gl_rom_n_1430, ZN => gl_rom_n_1467);
  gl_rom_g34951 : ND4D0BWP7T port map(A1 => gl_rom_n_1359, A2 => gl_rom_n_1429, A3 => gl_rom_n_1360, A4 => gl_rom_n_1356, ZN => gl_rom_n_1466);
  gl_rom_g34952 : ND4D0BWP7T port map(A1 => gl_rom_n_1426, A2 => gl_rom_n_1344, A3 => gl_rom_n_1347, A4 => gl_rom_n_1355, ZN => gl_rom_n_1465);
  gl_rom_g34953 : ND4D0BWP7T port map(A1 => gl_rom_n_1425, A2 => gl_rom_n_1346, A3 => gl_rom_n_1343, A4 => gl_rom_n_1348, ZN => gl_rom_n_1464);
  gl_rom_g34954 : ND4D0BWP7T port map(A1 => gl_rom_n_1446, A2 => gl_rom_n_1414, A3 => gl_rom_n_1408, A4 => gl_rom_n_1405, ZN => gl_rom_n_1463);
  gl_rom_g34955 : ND4D0BWP7T port map(A1 => gl_rom_n_1413, A2 => gl_rom_n_1415, A3 => gl_rom_n_1410, A4 => gl_rom_n_1412, ZN => gl_rom_n_1462);
  gl_rom_g34956 : ND4D0BWP7T port map(A1 => gl_rom_n_1330, A2 => gl_rom_n_1419, A3 => gl_rom_n_1327, A4 => gl_rom_n_1325, ZN => gl_rom_n_1461);
  gl_rom_g34957 : ND4D0BWP7T port map(A1 => gl_rom_n_1329, A2 => gl_rom_n_1320, A3 => gl_rom_n_1418, A4 => gl_rom_n_1326, ZN => gl_rom_n_1460);
  gl_rom_g34958 : ND4D0BWP7T port map(A1 => gl_rom_n_1324, A2 => gl_rom_n_1323, A3 => gl_rom_n_1319, A4 => gl_rom_n_1417, ZN => gl_rom_n_1459);
  gl_rom_g34959 : ND4D0BWP7T port map(A1 => gl_rom_n_1373, A2 => gl_rom_n_1322, A3 => gl_rom_n_1441, A4 => gl_rom_n_1351, ZN => gl_rom_n_1458);
  gl_rom_g34960 : ND4D0BWP7T port map(A1 => gl_rom_n_1411, A2 => gl_rom_n_1444, A3 => gl_rom_n_1399, A4 => gl_rom_n_1393, ZN => gl_rom_n_1457);
  gl_rom_g34961 : ND4D0BWP7T port map(A1 => gl_rom_n_1387, A2 => gl_rom_n_1388, A3 => gl_rom_n_1439, A4 => gl_rom_n_1390, ZN => gl_rom_n_1456);
  gl_rom_g34962 : ND4D0BWP7T port map(A1 => gl_rom_n_1389, A2 => gl_rom_n_1384, A3 => gl_rom_n_1380, A4 => gl_rom_n_1438, ZN => gl_rom_n_1455);
  gl_rom_g34963 : ND4D0BWP7T port map(A1 => gl_rom_n_1423, A2 => gl_rom_n_1361, A3 => gl_rom_n_1402, A4 => gl_rom_n_1353, ZN => gl_rom_n_1454);
  gl_rom_g34964 : ND4D0BWP7T port map(A1 => gl_rom_n_1432, A2 => gl_rom_n_1364, A3 => gl_rom_n_1367, A4 => gl_rom_n_1362, ZN => gl_rom_n_1453);
  gl_rom_g34965 : ND4D0BWP7T port map(A1 => gl_rom_n_1431, A2 => gl_rom_n_1358, A3 => gl_rom_n_1345, A4 => gl_rom_n_1382, ZN => gl_rom_n_1452);
  gl_rom_g34966 : ND4D0BWP7T port map(A1 => gl_rom_n_1354, A2 => gl_rom_n_1352, A3 => gl_rom_n_1349, A4 => gl_rom_n_1428, ZN => gl_rom_n_1451);
  gl_rom_g34967 : ND4D0BWP7T port map(A1 => gl_rom_n_1422, A2 => gl_rom_n_1333, A3 => gl_rom_n_1328, A4 => gl_rom_n_1321, ZN => gl_rom_n_1450);
  gl_rom_g34968 : ND4D0BWP7T port map(A1 => gl_rom_n_1336, A2 => gl_rom_n_1421, A3 => gl_rom_n_1331, A4 => gl_rom_n_1335, ZN => gl_rom_n_1449);
  gl_rom_g34969 : ND4D0BWP7T port map(A1 => gl_rom_n_1334, A2 => gl_rom_n_1416, A3 => gl_rom_n_1406, A4 => gl_rom_n_1395, ZN => gl_rom_n_1448);
  gl_rom_g34970 : ND4D0BWP7T port map(A1 => gl_rom_n_1338, A2 => gl_rom_n_1420, A3 => gl_rom_n_1332, A4 => gl_rom_n_1339, ZN => gl_rom_n_1447);
  gl_rom_g34971 : AOI22D0BWP7T port map(A1 => gl_rom_n_1312, A2 => gl_rom_n_26, B1 => gl_rom_n_1314, B2 => gl_rom_n_27, ZN => gl_rom_n_1446);
  gl_rom_g34972 : AOI22D0BWP7T port map(A1 => gl_rom_n_1295, A2 => gl_rom_n_25, B1 => gl_rom_n_1297, B2 => gl_rom_n_28, ZN => gl_rom_n_1445);
  gl_rom_g34973 : AOI22D0BWP7T port map(A1 => gl_rom_n_1284, A2 => gl_rom_n_25, B1 => gl_rom_n_1290, B2 => gl_rom_n_28, ZN => gl_rom_n_1444);
  gl_rom_g34974 : AOI22D0BWP7T port map(A1 => gl_rom_n_1282, A2 => gl_rom_n_25, B1 => gl_rom_n_1285, B2 => gl_rom_n_28, ZN => gl_rom_n_1443);
  gl_rom_g34975 : AOI22D0BWP7T port map(A1 => gl_rom_n_1273, A2 => gl_rom_n_25, B1 => gl_rom_n_1276, B2 => gl_rom_n_28, ZN => gl_rom_n_1442);
  gl_rom_g34976 : AOI22D0BWP7T port map(A1 => gl_rom_n_1231, A2 => gl_rom_n_25, B1 => gl_rom_n_1264, B2 => gl_rom_n_28, ZN => gl_rom_n_1441);
  gl_rom_g34977 : AOI22D0BWP7T port map(A1 => gl_rom_n_1268, A2 => gl_rom_n_25, B1 => gl_rom_n_1270, B2 => gl_rom_n_28, ZN => gl_rom_n_1440);
  gl_rom_g34978 : AOI22D0BWP7T port map(A1 => gl_rom_n_1254, A2 => gl_rom_n_25, B1 => gl_rom_n_1255, B2 => gl_rom_n_28, ZN => gl_rom_n_1439);
  gl_rom_g34979 : AOI22D0BWP7T port map(A1 => gl_rom_n_1240, A2 => gl_rom_n_25, B1 => gl_rom_n_1244, B2 => gl_rom_n_28, ZN => gl_rom_n_1438);
  gl_rom_g34980 : AOI22D0BWP7T port map(A1 => gl_rom_n_1232, A2 => gl_rom_n_25, B1 => gl_rom_n_1233, B2 => gl_rom_n_28, ZN => gl_rom_n_1437);
  gl_rom_g34981 : AOI22D0BWP7T port map(A1 => gl_rom_n_1219, A2 => gl_rom_n_25, B1 => gl_rom_n_1222, B2 => gl_rom_n_28, ZN => gl_rom_n_1436);
  gl_rom_g34982 : AOI22D0BWP7T port map(A1 => gl_rom_n_1207, A2 => gl_rom_n_25, B1 => gl_rom_n_1212, B2 => gl_rom_n_28, ZN => gl_rom_n_1435);
  gl_rom_g34983 : AOI22D0BWP7T port map(A1 => gl_rom_n_1203, A2 => gl_rom_n_25, B1 => gl_rom_n_1205, B2 => gl_rom_n_28, ZN => gl_rom_n_1434);
  gl_rom_g34984 : AOI22D0BWP7T port map(A1 => gl_rom_n_1204, A2 => gl_rom_n_25, B1 => gl_rom_n_1206, B2 => gl_rom_n_28, ZN => gl_rom_n_1433);
  gl_rom_g34985 : AOI22D0BWP7T port map(A1 => gl_rom_n_1187, A2 => gl_rom_n_25, B1 => gl_rom_n_1189, B2 => gl_rom_n_28, ZN => gl_rom_n_1432);
  gl_rom_g34986 : AOI22D0BWP7T port map(A1 => gl_rom_n_1172, A2 => gl_rom_n_25, B1 => gl_rom_n_1180, B2 => gl_rom_n_28, ZN => gl_rom_n_1431);
  gl_rom_g34987 : AOI22D0BWP7T port map(A1 => gl_rom_n_1169, A2 => gl_rom_n_25, B1 => gl_rom_n_1173, B2 => gl_rom_n_28, ZN => gl_rom_n_1430);
  gl_rom_g34988 : AOI22D0BWP7T port map(A1 => gl_rom_n_1167, A2 => gl_rom_n_25, B1 => gl_rom_n_1168, B2 => gl_rom_n_28, ZN => gl_rom_n_1429);
  gl_rom_g34989 : AOI22D0BWP7T port map(A1 => gl_rom_n_1159, A2 => gl_rom_n_25, B1 => gl_rom_n_1160, B2 => gl_rom_n_28, ZN => gl_rom_n_1428);
  gl_rom_g34990 : AOI22D0BWP7T port map(A1 => gl_rom_n_1151, A2 => gl_rom_n_25, B1 => gl_rom_n_1165, B2 => gl_rom_n_28, ZN => gl_rom_n_1427);
  gl_rom_g34991 : AOI22D0BWP7T port map(A1 => gl_rom_n_1146, A2 => gl_rom_n_25, B1 => gl_rom_n_1149, B2 => gl_rom_n_28, ZN => gl_rom_n_1426);
  gl_rom_g34992 : AOI22D0BWP7T port map(A1 => gl_rom_n_1140, A2 => gl_rom_n_25, B1 => gl_rom_n_1142, B2 => gl_rom_n_28, ZN => gl_rom_n_1425);
  gl_rom_g34993 : AOI22D0BWP7T port map(A1 => gl_rom_n_1119, A2 => gl_rom_n_25, B1 => gl_rom_n_1120, B2 => gl_rom_n_28, ZN => gl_rom_n_1424);
  gl_rom_g34994 : AOI22D0BWP7T port map(A1 => gl_rom_n_1191, A2 => gl_rom_n_25, B1 => gl_rom_n_1085, B2 => gl_rom_n_28, ZN => gl_rom_n_1423);
  gl_rom_g34995 : AOI22D0BWP7T port map(A1 => gl_rom_n_1109, A2 => gl_rom_n_25, B1 => gl_rom_n_1115, B2 => gl_rom_n_28, ZN => gl_rom_n_1422);
  gl_rom_g34996 : AOI22D0BWP7T port map(A1 => gl_rom_n_1106, A2 => gl_rom_n_25, B1 => gl_rom_n_1110, B2 => gl_rom_n_28, ZN => gl_rom_n_1421);
  gl_rom_g34997 : AOI22D0BWP7T port map(A1 => gl_rom_n_1105, A2 => gl_rom_n_25, B1 => gl_rom_n_1107, B2 => gl_rom_n_28, ZN => gl_rom_n_1420);
  gl_rom_g34998 : AOI22D0BWP7T port map(A1 => gl_rom_n_1091, A2 => gl_rom_n_25, B1 => gl_rom_n_1093, B2 => gl_rom_n_28, ZN => gl_rom_n_1419);
  gl_rom_g34999 : AOI22D0BWP7T port map(A1 => gl_rom_n_1073, A2 => gl_rom_n_25, B1 => gl_rom_n_1075, B2 => gl_rom_n_28, ZN => gl_rom_n_1418);
  gl_rom_g35000 : AOI22D0BWP7T port map(A1 => gl_rom_n_1071, A2 => gl_rom_n_25, B1 => gl_rom_n_1072, B2 => gl_rom_n_28, ZN => gl_rom_n_1417);
  gl_rom_g35001 : AOI22D0BWP7T port map(A1 => gl_rom_n_1308, A2 => gl_rom_n_25, B1 => gl_rom_n_1067, B2 => gl_rom_n_28, ZN => gl_rom_n_1416);
  gl_rom_g35002 : AOI22D0BWP7T port map(A1 => gl_rom_n_1317, A2 => gl_rom_n_25, B1 => gl_rom_n_1190, B2 => gl_rom_n_28, ZN => gl_rom_n_1415);
  gl_rom_g35003 : AOI22D0BWP7T port map(A1 => gl_rom_n_1304, A2 => gl_rom_n_25, B1 => gl_rom_n_1307, B2 => gl_rom_n_28, ZN => gl_rom_n_1414);
  gl_rom_g35004 : AOI22D0BWP7T port map(A1 => gl_rom_n_1313, A2 => gl_rom_n_23, B1 => gl_rom_n_1315, B2 => gl_rom_n_30, ZN => gl_rom_n_1413);
  gl_rom_g35005 : AOI22D0BWP7T port map(A1 => gl_rom_n_1310, A2 => gl_rom_n_26, B1 => gl_rom_n_1311, B2 => gl_rom_n_27, ZN => gl_rom_n_1412);
  gl_rom_g35006 : AOI22D0BWP7T port map(A1 => gl_rom_n_1300, A2 => gl_rom_n_23, B1 => gl_rom_n_1306, B2 => gl_rom_n_30, ZN => gl_rom_n_1411);
  gl_rom_g35007 : AOI22D0BWP7T port map(A1 => gl_rom_n_1305, A2 => gl_rom_n_24, B1 => gl_rom_n_1309, B2 => gl_rom_n_29, ZN => gl_rom_n_1410);
  gl_rom_g35008 : AOI22D0BWP7T port map(A1 => gl_rom_n_1302, A2 => gl_rom_n_26, B1 => gl_rom_n_1303, B2 => gl_rom_n_27, ZN => gl_rom_n_1409);
  gl_rom_g35009 : AOI22D0BWP7T port map(A1 => gl_rom_n_1296, A2 => gl_rom_n_23, B1 => gl_rom_n_1299, B2 => gl_rom_n_30, ZN => gl_rom_n_1408);
  gl_rom_g35010 : AOI22D0BWP7T port map(A1 => gl_rom_n_1298, A2 => gl_rom_n_23, B1 => gl_rom_n_1301, B2 => gl_rom_n_30, ZN => gl_rom_n_1407);
  gl_rom_g35011 : AOI22D0BWP7T port map(A1 => gl_rom_n_1277, A2 => gl_rom_n_26, B1 => gl_rom_n_1291, B2 => gl_rom_n_27, ZN => gl_rom_n_1406);
  gl_rom_g35012 : AOI22D0BWP7T port map(A1 => gl_rom_n_1288, A2 => gl_rom_n_24, B1 => gl_rom_n_1292, B2 => gl_rom_n_29, ZN => gl_rom_n_1405);
  gl_rom_g35013 : AOI22D0BWP7T port map(A1 => gl_rom_n_1289, A2 => gl_rom_n_24, B1 => gl_rom_n_1293, B2 => gl_rom_n_29, ZN => gl_rom_n_1404);
  gl_rom_g35014 : AOI22D0BWP7T port map(A1 => gl_rom_n_1286, A2 => gl_rom_n_26, B1 => gl_rom_n_1287, B2 => gl_rom_n_27, ZN => gl_rom_n_1403);
  gl_rom_g35015 : AOI22D0BWP7T port map(A1 => gl_rom_n_1200, A2 => gl_rom_n_26, B1 => gl_rom_n_1262, B2 => gl_rom_n_27, ZN => gl_rom_n_1402);
  gl_rom_g35016 : AOI22D0BWP7T port map(A1 => gl_rom_n_1281, A2 => gl_rom_n_26, B1 => gl_rom_n_1283, B2 => gl_rom_n_27, ZN => gl_rom_n_1401);
  gl_rom_g35017 : AOI22D0BWP7T port map(A1 => gl_rom_n_1279, A2 => gl_rom_n_23, B1 => gl_rom_n_1280, B2 => gl_rom_n_30, ZN => gl_rom_n_1400);
  gl_rom_g35018 : AOI22D0BWP7T port map(A1 => gl_rom_n_1267, A2 => gl_rom_n_26, B1 => gl_rom_n_1275, B2 => gl_rom_n_27, ZN => gl_rom_n_1399);
  gl_rom_g35019 : AOI22D0BWP7T port map(A1 => gl_rom_n_1274, A2 => gl_rom_n_24, B1 => gl_rom_n_1278, B2 => gl_rom_n_29, ZN => gl_rom_n_1398);
  gl_rom_g35020 : AOI22D0BWP7T port map(A1 => gl_rom_n_1271, A2 => gl_rom_n_26, B1 => gl_rom_n_1272, B2 => gl_rom_n_27, ZN => gl_rom_n_1397);
  gl_rom_g35021 : AOI22D0BWP7T port map(A1 => gl_rom_n_1265, A2 => gl_rom_n_23, B1 => gl_rom_n_1269, B2 => gl_rom_n_30, ZN => gl_rom_n_1396);
  gl_rom_g35022 : AOI22D0BWP7T port map(A1 => gl_rom_n_1245, A2 => gl_rom_n_24, B1 => gl_rom_n_1261, B2 => gl_rom_n_29, ZN => gl_rom_n_1395);
  gl_rom_g35023 : AOI22D0BWP7T port map(A1 => gl_rom_n_1263, A2 => gl_rom_n_23, B1 => gl_rom_n_1266, B2 => gl_rom_n_30, ZN => gl_rom_n_1394);
  gl_rom_g35024 : AOI22D0BWP7T port map(A1 => gl_rom_n_1253, A2 => gl_rom_n_24, B1 => gl_rom_n_1259, B2 => gl_rom_n_29, ZN => gl_rom_n_1393);
  gl_rom_g35025 : AOI22D0BWP7T port map(A1 => gl_rom_n_1256, A2 => gl_rom_n_24, B1 => gl_rom_n_1258, B2 => gl_rom_n_29, ZN => gl_rom_n_1392);
  gl_rom_g35026 : AOI22D0BWP7T port map(A1 => gl_rom_n_1257, A2 => gl_rom_n_24, B1 => gl_rom_n_1260, B2 => gl_rom_n_29, ZN => gl_rom_n_1391);
  gl_rom_g35027 : AOI22D0BWP7T port map(A1 => gl_rom_n_1250, A2 => gl_rom_n_23, B1 => gl_rom_n_1252, B2 => gl_rom_n_30, ZN => gl_rom_n_1390);
  gl_rom_g35028 : AOI22D0BWP7T port map(A1 => gl_rom_n_1249, A2 => gl_rom_n_23, B1 => gl_rom_n_1251, B2 => gl_rom_n_30, ZN => gl_rom_n_1389);
  gl_rom_g35029 : AOI22D0BWP7T port map(A1 => gl_rom_n_1247, A2 => gl_rom_n_26, B1 => gl_rom_n_1248, B2 => gl_rom_n_27, ZN => gl_rom_n_1388);
  gl_rom_g35030 : AOI22D0BWP7T port map(A1 => gl_rom_n_1242, A2 => gl_rom_n_24, B1 => gl_rom_n_1246, B2 => gl_rom_n_29, ZN => gl_rom_n_1387);
  gl_rom_g35031 : AOI22D0BWP7T port map(A1 => gl_rom_n_1238, A2 => gl_rom_n_26, B1 => gl_rom_n_1243, B2 => gl_rom_n_27, ZN => gl_rom_n_1386);
  gl_rom_g35032 : AOI22D0BWP7T port map(A1 => gl_rom_n_1239, A2 => gl_rom_n_26, B1 => gl_rom_n_1241, B2 => gl_rom_n_27, ZN => gl_rom_n_1385);
  gl_rom_g35033 : AOI22D0BWP7T port map(A1 => gl_rom_n_1234, A2 => gl_rom_n_26, B1 => gl_rom_n_1236, B2 => gl_rom_n_27, ZN => gl_rom_n_1384);
  gl_rom_g35034 : AOI22D0BWP7T port map(A1 => gl_rom_n_1235, A2 => gl_rom_n_23, B1 => gl_rom_n_1237, B2 => gl_rom_n_30, ZN => gl_rom_n_1383);
  gl_rom_g35035 : AOI22D0BWP7T port map(A1 => gl_rom_n_1143, A2 => gl_rom_n_26, B1 => gl_rom_n_1148, B2 => gl_rom_n_27, ZN => gl_rom_n_1382);
  gl_rom_g35036 : AOI22D0BWP7T port map(A1 => gl_rom_n_1220, A2 => gl_rom_n_23, B1 => gl_rom_n_1227, B2 => gl_rom_n_30, ZN => gl_rom_n_1381);
  gl_rom_g35037 : AOI22D0BWP7T port map(A1 => gl_rom_n_1226, A2 => gl_rom_n_24, B1 => gl_rom_n_1229, B2 => gl_rom_n_29, ZN => gl_rom_n_1380);
  gl_rom_g35038 : AOI22D0BWP7T port map(A1 => gl_rom_n_1228, A2 => gl_rom_n_24, B1 => gl_rom_n_1230, B2 => gl_rom_n_29, ZN => gl_rom_n_1379);
  gl_rom_g35039 : AOI22D0BWP7T port map(A1 => gl_rom_n_1224, A2 => gl_rom_n_26, B1 => gl_rom_n_1225, B2 => gl_rom_n_27, ZN => gl_rom_n_1378);
  gl_rom_g35040 : AOI22D0BWP7T port map(A1 => gl_rom_n_1218, A2 => gl_rom_n_26, B1 => gl_rom_n_1221, B2 => gl_rom_n_27, ZN => gl_rom_n_1377);
  gl_rom_g35041 : AOI22D0BWP7T port map(A1 => gl_rom_n_1209, A2 => gl_rom_n_23, B1 => gl_rom_n_1213, B2 => gl_rom_n_30, ZN => gl_rom_n_1376);
  gl_rom_g35042 : AOI22D0BWP7T port map(A1 => gl_rom_n_1216, A2 => gl_rom_n_23, B1 => gl_rom_n_1217, B2 => gl_rom_n_30, ZN => gl_rom_n_1375);
  gl_rom_g35043 : AOI22D0BWP7T port map(A1 => gl_rom_n_1211, A2 => gl_rom_n_24, B1 => gl_rom_n_1215, B2 => gl_rom_n_29, ZN => gl_rom_n_1374);
  gl_rom_g35044 : AOI22D0BWP7T port map(A1 => gl_rom_n_1170, A2 => gl_rom_n_23, B1 => gl_rom_n_1199, B2 => gl_rom_n_30, ZN => gl_rom_n_1373);
  gl_rom_g35045 : AOI22D0BWP7T port map(A1 => gl_rom_n_1208, A2 => gl_rom_n_26, B1 => gl_rom_n_1210, B2 => gl_rom_n_27, ZN => gl_rom_n_1372);
  gl_rom_g35046 : AOI22D0BWP7T port map(A1 => gl_rom_n_1183, A2 => gl_rom_n_23, B1 => gl_rom_n_1197, B2 => gl_rom_n_30, ZN => gl_rom_n_1371);
  gl_rom_g35047 : AOI22D0BWP7T port map(A1 => gl_rom_n_1201, A2 => gl_rom_n_23, B1 => gl_rom_n_1202, B2 => gl_rom_n_30, ZN => gl_rom_n_1370);
  gl_rom_g35048 : AOI22D0BWP7T port map(A1 => gl_rom_n_1194, A2 => gl_rom_n_24, B1 => gl_rom_n_1198, B2 => gl_rom_n_29, ZN => gl_rom_n_1369);
  gl_rom_g35049 : AOI22D0BWP7T port map(A1 => gl_rom_n_1193, A2 => gl_rom_n_24, B1 => gl_rom_n_1196, B2 => gl_rom_n_29, ZN => gl_rom_n_1368);
  gl_rom_g35050 : AOI22D0BWP7T port map(A1 => gl_rom_n_1318, A2 => gl_rom_n_23, B1 => gl_rom_n_1192, B2 => gl_rom_n_30, ZN => gl_rom_n_1367);
  gl_rom_g35051 : AOI22D0BWP7T port map(A1 => gl_rom_n_1063, A2 => gl_rom_n_24, B1 => gl_rom_n_1195, B2 => gl_rom_n_29, ZN => gl_rom_n_1366);
  gl_rom_g35052 : AOI22D0BWP7T port map(A1 => gl_rom_n_1185, A2 => gl_rom_n_26, B1 => gl_rom_n_1188, B2 => gl_rom_n_27, ZN => gl_rom_n_1365);
  gl_rom_g35053 : AOI22D0BWP7T port map(A1 => gl_rom_n_1184, A2 => gl_rom_n_26, B1 => gl_rom_n_1186, B2 => gl_rom_n_27, ZN => gl_rom_n_1364);
  gl_rom_g35054 : AOI22D0BWP7T port map(A1 => gl_rom_n_1177, A2 => gl_rom_n_23, B1 => gl_rom_n_1181, B2 => gl_rom_n_30, ZN => gl_rom_n_1363);
  gl_rom_g35055 : AOI22D0BWP7T port map(A1 => gl_rom_n_1179, A2 => gl_rom_n_24, B1 => gl_rom_n_1182, B2 => gl_rom_n_29, ZN => gl_rom_n_1362);
  gl_rom_g35056 : AOI22D0BWP7T port map(A1 => gl_rom_n_1087, A2 => gl_rom_n_23, B1 => gl_rom_n_1178, B2 => gl_rom_n_30, ZN => gl_rom_n_1361);
  gl_rom_g35057 : AOI22D0BWP7T port map(A1 => gl_rom_n_1175, A2 => gl_rom_n_26, B1 => gl_rom_n_1176, B2 => gl_rom_n_27, ZN => gl_rom_n_1360);
  gl_rom_g35058 : AOI22D0BWP7T port map(A1 => gl_rom_n_1171, A2 => gl_rom_n_23, B1 => gl_rom_n_1174, B2 => gl_rom_n_30, ZN => gl_rom_n_1359);
  gl_rom_g35059 : AOI22D0BWP7T port map(A1 => gl_rom_n_1156, A2 => gl_rom_n_23, B1 => gl_rom_n_1163, B2 => gl_rom_n_30, ZN => gl_rom_n_1358);
  gl_rom_g35060 : AOI22D0BWP7T port map(A1 => gl_rom_n_1161, A2 => gl_rom_n_24, B1 => gl_rom_n_1164, B2 => gl_rom_n_29, ZN => gl_rom_n_1357);
  gl_rom_g35061 : AOI22D0BWP7T port map(A1 => gl_rom_n_1162, A2 => gl_rom_n_24, B1 => gl_rom_n_1166, B2 => gl_rom_n_29, ZN => gl_rom_n_1356);
  gl_rom_g35062 : AOI22D0BWP7T port map(A1 => gl_rom_n_1153, A2 => gl_rom_n_26, B1 => gl_rom_n_1157, B2 => gl_rom_n_27, ZN => gl_rom_n_1355);
  gl_rom_g35063 : AOI22D0BWP7T port map(A1 => gl_rom_n_1155, A2 => gl_rom_n_23, B1 => gl_rom_n_1158, B2 => gl_rom_n_30, ZN => gl_rom_n_1354);
  gl_rom_g35064 : AOI22D0BWP7T port map(A1 => gl_rom_n_1108, A2 => gl_rom_n_24, B1 => gl_rom_n_1139, B2 => gl_rom_n_29, ZN => gl_rom_n_1353);
  gl_rom_g35065 : AOI22D0BWP7T port map(A1 => gl_rom_n_1152, A2 => gl_rom_n_26, B1 => gl_rom_n_1154, B2 => gl_rom_n_27, ZN => gl_rom_n_1352);
  gl_rom_g35066 : AOI22D0BWP7T port map(A1 => gl_rom_n_1118, A2 => gl_rom_n_24, B1 => gl_rom_n_1135, B2 => gl_rom_n_29, ZN => gl_rom_n_1351);
  gl_rom_g35067 : AOI22D0BWP7T port map(A1 => gl_rom_n_1214, A2 => gl_rom_n_26, B1 => gl_rom_n_1223, B2 => gl_rom_n_27, ZN => gl_rom_n_1350);
  gl_rom_g35068 : AOI22D0BWP7T port map(A1 => gl_rom_n_1147, A2 => gl_rom_n_24, B1 => gl_rom_n_1150, B2 => gl_rom_n_29, ZN => gl_rom_n_1349);
  gl_rom_g35069 : AOI22D0BWP7T port map(A1 => gl_rom_n_1144, A2 => gl_rom_n_26, B1 => gl_rom_n_1145, B2 => gl_rom_n_27, ZN => gl_rom_n_1348);
  gl_rom_g35070 : AOI22D0BWP7T port map(A1 => gl_rom_n_1138, A2 => gl_rom_n_23, B1 => gl_rom_n_1141, B2 => gl_rom_n_30, ZN => gl_rom_n_1347);
  gl_rom_g35071 : AOI22D0BWP7T port map(A1 => gl_rom_n_1136, A2 => gl_rom_n_23, B1 => gl_rom_n_1137, B2 => gl_rom_n_30, ZN => gl_rom_n_1346);
  gl_rom_g35072 : AOI22D0BWP7T port map(A1 => gl_rom_n_1128, A2 => gl_rom_n_24, B1 => gl_rom_n_1131, B2 => gl_rom_n_29, ZN => gl_rom_n_1345);
  gl_rom_g35073 : AOI22D0BWP7T port map(A1 => gl_rom_n_1129, A2 => gl_rom_n_24, B1 => gl_rom_n_1132, B2 => gl_rom_n_29, ZN => gl_rom_n_1344);
  gl_rom_g35074 : AOI22D0BWP7T port map(A1 => gl_rom_n_1130, A2 => gl_rom_n_24, B1 => gl_rom_n_1134, B2 => gl_rom_n_29, ZN => gl_rom_n_1343);
  gl_rom_g35075 : AOI22D0BWP7T port map(A1 => gl_rom_n_1126, A2 => gl_rom_n_26, B1 => gl_rom_n_1127, B2 => gl_rom_n_27, ZN => gl_rom_n_1342);
  gl_rom_g35076 : AOI22D0BWP7T port map(A1 => gl_rom_n_1125, A2 => gl_rom_n_24, B1 => gl_rom_n_1133, B2 => gl_rom_n_29, ZN => gl_rom_n_1341);
  gl_rom_g35077 : AOI22D0BWP7T port map(A1 => gl_rom_n_1122, A2 => gl_rom_n_23, B1 => gl_rom_n_1124, B2 => gl_rom_n_30, ZN => gl_rom_n_1340);
  gl_rom_g35078 : AOI22D0BWP7T port map(A1 => gl_rom_n_1121, A2 => gl_rom_n_26, B1 => gl_rom_n_1123, B2 => gl_rom_n_27, ZN => gl_rom_n_1339);
  gl_rom_g35079 : AOI22D0BWP7T port map(A1 => gl_rom_n_1113, A2 => gl_rom_n_23, B1 => gl_rom_n_1116, B2 => gl_rom_n_30, ZN => gl_rom_n_1338);
  gl_rom_g35080 : AOI22D0BWP7T port map(A1 => gl_rom_n_1114, A2 => gl_rom_n_24, B1 => gl_rom_n_1117, B2 => gl_rom_n_29, ZN => gl_rom_n_1337);
  gl_rom_g35081 : AOI22D0BWP7T port map(A1 => gl_rom_n_1111, A2 => gl_rom_n_23, B1 => gl_rom_n_1112, B2 => gl_rom_n_30, ZN => gl_rom_n_1336);
  gl_rom_g35082 : AOI22D0BWP7T port map(A1 => gl_rom_n_1103, A2 => gl_rom_n_26, B1 => gl_rom_n_1104, B2 => gl_rom_n_27, ZN => gl_rom_n_1335);
  gl_rom_g35083 : AOI22D0BWP7T port map(A1 => gl_rom_n_1084, A2 => gl_rom_n_23, B1 => gl_rom_n_1099, B2 => gl_rom_n_30, ZN => gl_rom_n_1334);
  gl_rom_g35084 : AOI22D0BWP7T port map(A1 => gl_rom_n_1094, A2 => gl_rom_n_23, B1 => gl_rom_n_1101, B2 => gl_rom_n_30, ZN => gl_rom_n_1333);
  gl_rom_g35085 : AOI22D0BWP7T port map(A1 => gl_rom_n_1096, A2 => gl_rom_n_24, B1 => gl_rom_n_1100, B2 => gl_rom_n_29, ZN => gl_rom_n_1332);
  gl_rom_g35086 : AOI22D0BWP7T port map(A1 => gl_rom_n_1098, A2 => gl_rom_n_24, B1 => gl_rom_n_1102, B2 => gl_rom_n_29, ZN => gl_rom_n_1331);
  gl_rom_g35087 : AOI22D0BWP7T port map(A1 => gl_rom_n_1095, A2 => gl_rom_n_26, B1 => gl_rom_n_1097, B2 => gl_rom_n_27, ZN => gl_rom_n_1330);
  gl_rom_g35088 : AOI22D0BWP7T port map(A1 => gl_rom_n_1090, A2 => gl_rom_n_26, B1 => gl_rom_n_1092, B2 => gl_rom_n_27, ZN => gl_rom_n_1329);
  gl_rom_g35089 : AOI22D0BWP7T port map(A1 => gl_rom_n_1076, A2 => gl_rom_n_26, B1 => gl_rom_n_1083, B2 => gl_rom_n_27, ZN => gl_rom_n_1328);
  gl_rom_g35090 : AOI22D0BWP7T port map(A1 => gl_rom_n_1088, A2 => gl_rom_n_23, B1 => gl_rom_n_1089, B2 => gl_rom_n_30, ZN => gl_rom_n_1327);
  gl_rom_g35091 : AOI22D0BWP7T port map(A1 => gl_rom_n_1080, A2 => gl_rom_n_23, B1 => gl_rom_n_1082, B2 => gl_rom_n_30, ZN => gl_rom_n_1326);
  gl_rom_g35092 : AOI22D0BWP7T port map(A1 => gl_rom_n_1081, A2 => gl_rom_n_24, B1 => gl_rom_n_1086, B2 => gl_rom_n_29, ZN => gl_rom_n_1325);
  gl_rom_g35093 : AOI22D0BWP7T port map(A1 => gl_rom_n_1078, A2 => gl_rom_n_26, B1 => gl_rom_n_1079, B2 => gl_rom_n_27, ZN => gl_rom_n_1324);
  gl_rom_g35094 : AOI22D0BWP7T port map(A1 => gl_rom_n_1074, A2 => gl_rom_n_23, B1 => gl_rom_n_1077, B2 => gl_rom_n_30, ZN => gl_rom_n_1323);
  gl_rom_g35095 : AOI22D0BWP7T port map(A1 => gl_rom_n_1294, A2 => gl_rom_n_26, B1 => gl_rom_n_1065, B2 => gl_rom_n_27, ZN => gl_rom_n_1322);
  gl_rom_g35096 : AOI22D0BWP7T port map(A1 => gl_rom_n_1316, A2 => gl_rom_n_24, B1 => gl_rom_n_1069, B2 => gl_rom_n_29, ZN => gl_rom_n_1321);
  gl_rom_g35097 : AOI22D0BWP7T port map(A1 => gl_rom_n_1064, A2 => gl_rom_n_24, B1 => gl_rom_n_1068, B2 => gl_rom_n_29, ZN => gl_rom_n_1320);
  gl_rom_g35098 : AOI22D0BWP7T port map(A1 => gl_rom_n_1066, A2 => gl_rom_n_24, B1 => gl_rom_n_1070, B2 => gl_rom_n_29, ZN => gl_rom_n_1319);
  gl_rom_g35099 : ND4D0BWP7T port map(A1 => gl_rom_n_546, A2 => gl_rom_n_294, A3 => gl_rom_n_549, A4 => gl_rom_n_547, ZN => gl_rom_n_1318);
  gl_rom_g35100 : ND4D0BWP7T port map(A1 => gl_rom_n_1056, A2 => gl_rom_n_1060, A3 => gl_rom_n_1059, A4 => gl_rom_n_1057, ZN => gl_rom_n_1317);
  gl_rom_g35101 : ND4D0BWP7T port map(A1 => gl_rom_n_1052, A2 => gl_rom_n_1036, A3 => gl_rom_n_1046, A4 => gl_rom_n_1033, ZN => gl_rom_n_1316);
  gl_rom_g35102 : ND4D0BWP7T port map(A1 => gl_rom_n_1047, A2 => gl_rom_n_1051, A3 => gl_rom_n_1050, A4 => gl_rom_n_1048, ZN => gl_rom_n_1315);
  gl_rom_g35103 : ND4D0BWP7T port map(A1 => gl_rom_n_1049, A2 => gl_rom_n_1041, A3 => gl_rom_n_1045, A4 => gl_rom_n_1039, ZN => gl_rom_n_1314);
  gl_rom_g35104 : ND4D0BWP7T port map(A1 => gl_rom_n_1043, A2 => gl_rom_n_1044, A3 => gl_rom_n_1040, A4 => gl_rom_n_1038, ZN => gl_rom_n_1313);
  gl_rom_g35105 : ND4D0BWP7T port map(A1 => gl_rom_n_1030, A2 => gl_rom_n_1034, A3 => gl_rom_n_1026, A4 => gl_rom_n_1025, ZN => gl_rom_n_1312);
  gl_rom_g35106 : ND4D0BWP7T port map(A1 => gl_rom_n_1032, A2 => gl_rom_n_1035, A3 => gl_rom_n_1037, A4 => gl_rom_n_1031, ZN => gl_rom_n_1311);
  gl_rom_g35107 : ND4D0BWP7T port map(A1 => gl_rom_n_1024, A2 => gl_rom_n_1027, A3 => gl_rom_n_1029, A4 => gl_rom_n_1023, ZN => gl_rom_n_1310);
  gl_rom_g35108 : ND4D0BWP7T port map(A1 => gl_rom_n_1018, A2 => gl_rom_n_1020, A3 => gl_rom_n_1022, A4 => gl_rom_n_1016, ZN => gl_rom_n_1309);
  gl_rom_g35109 : ND4D0BWP7T port map(A1 => gl_rom_n_990, A2 => gl_rom_n_1010, A3 => gl_rom_n_1017, A4 => gl_rom_n_982, ZN => gl_rom_n_1308);
  gl_rom_g35110 : ND4D0BWP7T port map(A1 => gl_rom_n_1019, A2 => gl_rom_n_1012, A3 => gl_rom_n_1015, A4 => gl_rom_n_1007, ZN => gl_rom_n_1307);
  gl_rom_g35111 : ND4D0BWP7T port map(A1 => gl_rom_n_1005, A2 => gl_rom_n_1014, A3 => gl_rom_n_1004, A4 => gl_rom_n_998, ZN => gl_rom_n_1306);
  gl_rom_g35112 : ND4D0BWP7T port map(A1 => gl_rom_n_1009, A2 => gl_rom_n_1011, A3 => gl_rom_n_1013, A4 => gl_rom_n_1008, ZN => gl_rom_n_1305);
  gl_rom_g35113 : ND4D0BWP7T port map(A1 => gl_rom_n_1002, A2 => gl_rom_n_996, A3 => gl_rom_n_1000, A4 => gl_rom_n_993, ZN => gl_rom_n_1304);
  gl_rom_g35114 : ND4D0BWP7T port map(A1 => gl_rom_n_999, A2 => gl_rom_n_1006, A3 => gl_rom_n_1003, A4 => gl_rom_n_1001, ZN => gl_rom_n_1303);
  gl_rom_g35115 : ND4D0BWP7T port map(A1 => gl_rom_n_992, A2 => gl_rom_n_997, A3 => gl_rom_n_995, A4 => gl_rom_n_994, ZN => gl_rom_n_1302);
  gl_rom_g35116 : ND4D0BWP7T port map(A1 => gl_rom_n_986, A2 => gl_rom_n_989, A3 => gl_rom_n_991, A4 => gl_rom_n_984, ZN => gl_rom_n_1301);
  gl_rom_g35117 : ND4D0BWP7T port map(A1 => gl_rom_n_970, A2 => gl_rom_n_975, A3 => gl_rom_n_985, A4 => gl_rom_n_965, ZN => gl_rom_n_1300);
  gl_rom_g35118 : ND4D0BWP7T port map(A1 => gl_rom_n_987, A2 => gl_rom_n_979, A3 => gl_rom_n_983, A4 => gl_rom_n_977, ZN => gl_rom_n_1299);
  gl_rom_g35119 : ND4D0BWP7T port map(A1 => gl_rom_n_980, A2 => gl_rom_n_981, A3 => gl_rom_n_978, A4 => gl_rom_n_976, ZN => gl_rom_n_1298);
  gl_rom_g35120 : ND4D0BWP7T port map(A1 => gl_rom_n_967, A2 => gl_rom_n_974, A3 => gl_rom_n_972, A4 => gl_rom_n_969, ZN => gl_rom_n_1297);
  gl_rom_g35121 : ND4D0BWP7T port map(A1 => gl_rom_n_971, A2 => gl_rom_n_964, A3 => gl_rom_n_968, A4 => gl_rom_n_962, ZN => gl_rom_n_1296);
  gl_rom_g35122 : ND4D0BWP7T port map(A1 => gl_rom_n_963, A2 => gl_rom_n_960, A3 => gl_rom_n_966, A4 => gl_rom_n_961, ZN => gl_rom_n_1295);
  gl_rom_g35123 : ND4D0BWP7T port map(A1 => gl_rom_n_952, A2 => gl_rom_n_902, A3 => gl_rom_n_925, A4 => gl_rom_n_865, ZN => gl_rom_n_1294);
  gl_rom_g35124 : ND4D0BWP7T port map(A1 => gl_rom_n_956, A2 => gl_rom_n_958, A3 => gl_rom_n_959, A4 => gl_rom_n_955, ZN => gl_rom_n_1293);
  gl_rom_g35125 : ND4D0BWP7T port map(A1 => gl_rom_n_946, A2 => gl_rom_n_957, A3 => gl_rom_n_954, A4 => gl_rom_n_949, ZN => gl_rom_n_1292);
  gl_rom_g35126 : ND4D0BWP7T port map(A1 => gl_rom_n_950, A2 => gl_rom_n_928, A3 => gl_rom_n_943, A4 => gl_rom_n_910, ZN => gl_rom_n_1291);
  gl_rom_g35127 : ND4D0BWP7T port map(A1 => gl_rom_n_933, A2 => gl_rom_n_953, A3 => gl_rom_n_947, A4 => gl_rom_n_939, ZN => gl_rom_n_1290);
  gl_rom_g35128 : ND4D0BWP7T port map(A1 => gl_rom_n_948, A2 => gl_rom_n_951, A3 => gl_rom_n_945, A4 => gl_rom_n_944, ZN => gl_rom_n_1289);
  gl_rom_g35129 : ND4D0BWP7T port map(A1 => gl_rom_n_941, A2 => gl_rom_n_935, A3 => gl_rom_n_936, A4 => gl_rom_n_931, ZN => gl_rom_n_1288);
  gl_rom_g35130 : ND4D0BWP7T port map(A1 => gl_rom_n_938, A2 => gl_rom_n_940, A3 => gl_rom_n_942, A4 => gl_rom_n_937, ZN => gl_rom_n_1287);
  gl_rom_g35131 : ND4D0BWP7T port map(A1 => gl_rom_n_930, A2 => gl_rom_n_932, A3 => gl_rom_n_934, A4 => gl_rom_n_929, ZN => gl_rom_n_1286);
  gl_rom_g35132 : ND4D0BWP7T port map(A1 => gl_rom_n_927, A2 => gl_rom_n_923, A3 => gl_rom_n_926, A4 => gl_rom_n_922, ZN => gl_rom_n_1285);
  gl_rom_g35133 : ND4D0BWP7T port map(A1 => gl_rom_n_917, A2 => gl_rom_n_901, A3 => gl_rom_n_919, A4 => gl_rom_n_909, ZN => gl_rom_n_1284);
  gl_rom_g35134 : ND4D0BWP7T port map(A1 => gl_rom_n_916, A2 => gl_rom_n_921, A3 => gl_rom_n_924, A4 => gl_rom_n_915, ZN => gl_rom_n_1283);
  gl_rom_g35135 : ND4D0BWP7T port map(A1 => gl_rom_n_914, A2 => gl_rom_n_918, A3 => gl_rom_n_920, A4 => gl_rom_n_913, ZN => gl_rom_n_1282);
  gl_rom_g35136 : ND4D0BWP7T port map(A1 => gl_rom_n_906, A2 => gl_rom_n_898, A3 => gl_rom_n_907, A4 => gl_rom_n_900, ZN => gl_rom_n_1281);
  gl_rom_g35137 : ND4D0BWP7T port map(A1 => gl_rom_n_908, A2 => gl_rom_n_904, A3 => gl_rom_n_912, A4 => gl_rom_n_905, ZN => gl_rom_n_1280);
  gl_rom_g35138 : ND4D0BWP7T port map(A1 => gl_rom_n_897, A2 => gl_rom_n_899, A3 => gl_rom_n_903, A4 => gl_rom_n_896, ZN => gl_rom_n_1279);
  gl_rom_g35139 : ND4D0BWP7T port map(A1 => gl_rom_n_891, A2 => gl_rom_n_894, A3 => gl_rom_n_895, A4 => gl_rom_n_889, ZN => gl_rom_n_1278);
  gl_rom_g35140 : ND4D0BWP7T port map(A1 => gl_rom_n_879, A2 => gl_rom_n_846, A3 => gl_rom_n_893, A4 => gl_rom_n_864, ZN => gl_rom_n_1277);
  gl_rom_g35141 : ND4D0BWP7T port map(A1 => gl_rom_n_892, A2 => gl_rom_n_885, A3 => gl_rom_n_890, A4 => gl_rom_n_880, ZN => gl_rom_n_1276);
  gl_rom_g35142 : ND4D0BWP7T port map(A1 => gl_rom_n_872, A2 => gl_rom_n_888, A3 => gl_rom_n_887, A4 => gl_rom_n_876, ZN => gl_rom_n_1275);
  gl_rom_g35143 : ND4D0BWP7T port map(A1 => gl_rom_n_884, A2 => gl_rom_n_886, A3 => gl_rom_n_883, A4 => gl_rom_n_882, ZN => gl_rom_n_1274);
  gl_rom_g35144 : ND4D0BWP7T port map(A1 => gl_rom_n_878, A2 => gl_rom_n_871, A3 => gl_rom_n_874, A4 => gl_rom_n_867, ZN => gl_rom_n_1273);
  gl_rom_g35145 : ND4D0BWP7T port map(A1 => gl_rom_n_873, A2 => gl_rom_n_881, A3 => gl_rom_n_877, A4 => gl_rom_n_875, ZN => gl_rom_n_1272);
  gl_rom_g35146 : ND4D0BWP7T port map(A1 => gl_rom_n_869, A2 => gl_rom_n_870, A3 => gl_rom_n_868, A4 => gl_rom_n_866, ZN => gl_rom_n_1271);
  gl_rom_g35147 : ND4D0BWP7T port map(A1 => gl_rom_n_857, A2 => gl_rom_n_860, A3 => gl_rom_n_863, A4 => gl_rom_n_855, ZN => gl_rom_n_1270);
  gl_rom_g35148 : ND4D0BWP7T port map(A1 => gl_rom_n_859, A2 => gl_rom_n_853, A3 => gl_rom_n_856, A4 => gl_rom_n_848, ZN => gl_rom_n_1269);
  gl_rom_g35149 : ND4D0BWP7T port map(A1 => gl_rom_n_850, A2 => gl_rom_n_852, A3 => gl_rom_n_854, A4 => gl_rom_n_849, ZN => gl_rom_n_1268);
  gl_rom_g35150 : ND4D0BWP7T port map(A1 => gl_rom_n_851, A2 => gl_rom_n_838, A3 => gl_rom_n_858, A4 => gl_rom_n_845, ZN => gl_rom_n_1267);
  gl_rom_g35151 : ND4D0BWP7T port map(A1 => gl_rom_n_841, A2 => gl_rom_n_843, A3 => gl_rom_n_847, A4 => gl_rom_n_840, ZN => gl_rom_n_1266);
  gl_rom_g35152 : ND4D0BWP7T port map(A1 => gl_rom_n_837, A2 => gl_rom_n_842, A3 => gl_rom_n_844, A4 => gl_rom_n_835, ZN => gl_rom_n_1265);
  gl_rom_g35153 : ND4D0BWP7T port map(A1 => gl_rom_n_798, A2 => gl_rom_n_742, A3 => gl_rom_n_824, A4 => gl_rom_n_768, ZN => gl_rom_n_1264);
  gl_rom_g35154 : ND4D0BWP7T port map(A1 => gl_rom_n_834, A2 => gl_rom_n_836, A3 => gl_rom_n_839, A4 => gl_rom_n_833, ZN => gl_rom_n_1263);
  gl_rom_g35155 : ND4D0BWP7T port map(A1 => gl_rom_n_816, A2 => gl_rom_n_861, A3 => gl_rom_n_743, A4 => gl_rom_n_706, ZN => gl_rom_n_1262);
  gl_rom_g35156 : ND4D0BWP7T port map(A1 => gl_rom_n_811, A2 => gl_rom_n_783, A3 => gl_rom_n_829, A4 => gl_rom_n_800, ZN => gl_rom_n_1261);
  gl_rom_g35157 : ND4D0BWP7T port map(A1 => gl_rom_n_828, A2 => gl_rom_n_831, A3 => gl_rom_n_832, A4 => gl_rom_n_826, ZN => gl_rom_n_1260);
  gl_rom_g35158 : ND4D0BWP7T port map(A1 => gl_rom_n_817, A2 => gl_rom_n_827, A3 => gl_rom_n_814, A4 => gl_rom_n_1062, ZN => gl_rom_n_1259);
  gl_rom_g35159 : ND4D0BWP7T port map(A1 => gl_rom_n_825, A2 => gl_rom_n_820, A3 => gl_rom_n_830, A4 => gl_rom_n_822, ZN => gl_rom_n_1258);
  gl_rom_g35160 : ND4D0BWP7T port map(A1 => gl_rom_n_819, A2 => gl_rom_n_821, A3 => gl_rom_n_823, A4 => gl_rom_n_818, ZN => gl_rom_n_1257);
  gl_rom_g35161 : ND4D0BWP7T port map(A1 => gl_rom_n_815, A2 => gl_rom_n_807, A3 => gl_rom_n_810, A4 => gl_rom_n_803, ZN => gl_rom_n_1256);
  gl_rom_g35162 : ND4D0BWP7T port map(A1 => gl_rom_n_812, A2 => gl_rom_n_813, A3 => gl_rom_n_809, A4 => gl_rom_n_808, ZN => gl_rom_n_1255);
  gl_rom_g35163 : ND4D0BWP7T port map(A1 => gl_rom_n_802, A2 => gl_rom_n_804, A3 => gl_rom_n_805, A4 => gl_rom_n_801, ZN => gl_rom_n_1254);
  gl_rom_g35164 : ND4D0BWP7T port map(A1 => gl_rom_n_791, A2 => gl_rom_n_797, A3 => gl_rom_n_782, A4 => gl_rom_n_779, ZN => gl_rom_n_1253);
  gl_rom_g35165 : ND4D0BWP7T port map(A1 => gl_rom_n_799, A2 => gl_rom_n_794, A3 => gl_rom_n_796, A4 => gl_rom_n_793, ZN => gl_rom_n_1252);
  gl_rom_g35166 : ND4D0BWP7T port map(A1 => gl_rom_n_785, A2 => gl_rom_n_795, A3 => gl_rom_n_792, A4 => gl_rom_n_788, ZN => gl_rom_n_1251);
  gl_rom_g35167 : ND4D0BWP7T port map(A1 => gl_rom_n_787, A2 => gl_rom_n_789, A3 => gl_rom_n_790, A4 => gl_rom_n_786, ZN => gl_rom_n_1250);
  gl_rom_g35168 : ND4D0BWP7T port map(A1 => gl_rom_n_770, A2 => gl_rom_n_781, A3 => gl_rom_n_777, A4 => gl_rom_n_774, ZN => gl_rom_n_1249);
  gl_rom_g35169 : ND4D0BWP7T port map(A1 => gl_rom_n_784, A2 => gl_rom_n_778, A3 => gl_rom_n_780, A4 => gl_rom_n_776, ZN => gl_rom_n_1248);
  gl_rom_g35170 : ND4D0BWP7T port map(A1 => gl_rom_n_771, A2 => gl_rom_n_773, A3 => gl_rom_n_775, A4 => gl_rom_n_769, ZN => gl_rom_n_1247);
  gl_rom_g35171 : ND4D0BWP7T port map(A1 => gl_rom_n_765, A2 => gl_rom_n_766, A3 => gl_rom_n_763, A4 => gl_rom_n_762, ZN => gl_rom_n_1246);
  gl_rom_g35172 : ND4D0BWP7T port map(A1 => gl_rom_n_752, A2 => gl_rom_n_726, A3 => gl_rom_n_767, A4 => gl_rom_n_735, ZN => gl_rom_n_1245);
  gl_rom_g35173 : ND4D0BWP7T port map(A1 => gl_rom_n_761, A2 => gl_rom_n_764, A3 => gl_rom_n_758, A4 => gl_rom_n_754, ZN => gl_rom_n_1244);
  gl_rom_g35174 : ND4D0BWP7T port map(A1 => gl_rom_n_744, A2 => gl_rom_n_751, A3 => gl_rom_n_760, A4 => gl_rom_n_732, ZN => gl_rom_n_1243);
  gl_rom_g35175 : ND4D0BWP7T port map(A1 => gl_rom_n_755, A2 => gl_rom_n_757, A3 => gl_rom_n_759, A4 => gl_rom_n_753, ZN => gl_rom_n_1242);
  gl_rom_g35176 : ND4D0BWP7T port map(A1 => gl_rom_n_750, A2 => gl_rom_n_746, A3 => gl_rom_n_748, A4 => gl_rom_n_745, ZN => gl_rom_n_1241);
  gl_rom_g35177 : ND4D0BWP7T port map(A1 => gl_rom_n_740, A2 => gl_rom_n_747, A3 => gl_rom_n_749, A4 => gl_rom_n_736, ZN => gl_rom_n_1240);
  gl_rom_g35178 : ND4D0BWP7T port map(A1 => gl_rom_n_739, A2 => gl_rom_n_741, A3 => gl_rom_n_738, A4 => gl_rom_n_737, ZN => gl_rom_n_1239);
  gl_rom_g35179 : ND4D0BWP7T port map(A1 => gl_rom_n_708, A2 => gl_rom_n_727, A3 => gl_rom_n_722, A4 => gl_rom_n_712, ZN => gl_rom_n_1238);
  gl_rom_g35180 : ND4D0BWP7T port map(A1 => gl_rom_n_733, A2 => gl_rom_n_734, A3 => gl_rom_n_730, A4 => gl_rom_n_728, ZN => gl_rom_n_1237);
  gl_rom_g35181 : ND4D0BWP7T port map(A1 => gl_rom_n_724, A2 => gl_rom_n_729, A3 => gl_rom_n_731, A4 => gl_rom_n_719, ZN => gl_rom_n_1236);
  gl_rom_g35182 : ND4D0BWP7T port map(A1 => gl_rom_n_721, A2 => gl_rom_n_723, A3 => gl_rom_n_725, A4 => gl_rom_n_720, ZN => gl_rom_n_1235);
  gl_rom_g35183 : ND4D0BWP7T port map(A1 => gl_rom_n_705, A2 => gl_rom_n_716, A3 => gl_rom_n_714, A4 => gl_rom_n_710, ZN => gl_rom_n_1234);
  gl_rom_g35184 : ND4D0BWP7T port map(A1 => gl_rom_n_715, A2 => gl_rom_n_717, A3 => gl_rom_n_718, A4 => gl_rom_n_713, ZN => gl_rom_n_1233);
  gl_rom_g35185 : ND4D0BWP7T port map(A1 => gl_rom_n_709, A2 => gl_rom_n_711, A3 => gl_rom_n_707, A4 => gl_rom_n_704, ZN => gl_rom_n_1232);
  gl_rom_g35186 : ND4D0BWP7T port map(A1 => gl_rom_n_703, A2 => gl_rom_n_639, A3 => gl_rom_n_698, A4 => gl_rom_n_636, ZN => gl_rom_n_1231);
  gl_rom_g35187 : ND4D0BWP7T port map(A1 => gl_rom_n_699, A2 => gl_rom_n_701, A3 => gl_rom_n_702, A4 => gl_rom_n_696, ZN => gl_rom_n_1230);
  gl_rom_g35188 : ND4D0BWP7T port map(A1 => gl_rom_n_688, A2 => gl_rom_n_700, A3 => gl_rom_n_697, A4 => gl_rom_n_691, ZN => gl_rom_n_1229);
  gl_rom_g35189 : ND4D0BWP7T port map(A1 => gl_rom_n_690, A2 => gl_rom_n_692, A3 => gl_rom_n_694, A4 => gl_rom_n_687, ZN => gl_rom_n_1228);
  gl_rom_g35190 : ND4D0BWP7T port map(A1 => gl_rom_n_695, A2 => gl_rom_n_683, A3 => gl_rom_n_689, A4 => gl_rom_n_672, ZN => gl_rom_n_1227);
  gl_rom_g35191 : ND4D0BWP7T port map(A1 => gl_rom_n_675, A2 => gl_rom_n_686, A3 => gl_rom_n_682, A4 => gl_rom_n_678, ZN => gl_rom_n_1226);
  gl_rom_g35192 : ND4D0BWP7T port map(A1 => gl_rom_n_680, A2 => gl_rom_n_685, A3 => gl_rom_n_684, A4 => gl_rom_n_681, ZN => gl_rom_n_1225);
  gl_rom_g35193 : ND4D0BWP7T port map(A1 => gl_rom_n_676, A2 => gl_rom_n_673, A3 => gl_rom_n_677, A4 => gl_rom_n_674, ZN => gl_rom_n_1224);
  gl_rom_g35194 : ND4D0BWP7T port map(A1 => gl_rom_n_693, A2 => gl_rom_n_669, A3 => gl_rom_n_679, A4 => gl_rom_n_652, ZN => gl_rom_n_1223);
  gl_rom_g35195 : ND4D0BWP7T port map(A1 => gl_rom_n_666, A2 => gl_rom_n_671, A3 => gl_rom_n_670, A4 => gl_rom_n_667, ZN => gl_rom_n_1222);
  gl_rom_g35196 : ND4D0BWP7T port map(A1 => gl_rom_n_660, A2 => gl_rom_n_664, A3 => gl_rom_n_668, A4 => gl_rom_n_657, ZN => gl_rom_n_1221);
  gl_rom_g35197 : ND4D0BWP7T port map(A1 => gl_rom_n_665, A2 => gl_rom_n_655, A3 => gl_rom_n_663, A4 => gl_rom_n_648, ZN => gl_rom_n_1220);
  gl_rom_g35198 : ND4D0BWP7T port map(A1 => gl_rom_n_659, A2 => gl_rom_n_661, A3 => gl_rom_n_662, A4 => gl_rom_n_658, ZN => gl_rom_n_1219);
  gl_rom_g35199 : ND4D0BWP7T port map(A1 => gl_rom_n_645, A2 => gl_rom_n_650, A3 => gl_rom_n_653, A4 => gl_rom_n_643, ZN => gl_rom_n_1218);
  gl_rom_g35200 : ND4D0BWP7T port map(A1 => gl_rom_n_654, A2 => gl_rom_n_656, A3 => gl_rom_n_651, A4 => gl_rom_n_649, ZN => gl_rom_n_1217);
  gl_rom_g35201 : ND4D0BWP7T port map(A1 => gl_rom_n_647, A2 => gl_rom_n_644, A3 => gl_rom_n_646, A4 => gl_rom_n_642, ZN => gl_rom_n_1216);
  gl_rom_g35202 : ND4D0BWP7T port map(A1 => gl_rom_n_638, A2 => gl_rom_n_640, A3 => gl_rom_n_635, A4 => gl_rom_n_634, ZN => gl_rom_n_1215);
  gl_rom_g35203 : ND4D0BWP7T port map(A1 => gl_rom_n_589, A2 => gl_rom_n_628, A3 => gl_rom_n_623, A4 => gl_rom_n_608, ZN => gl_rom_n_1214);
  gl_rom_g35204 : ND4D0BWP7T port map(A1 => gl_rom_n_627, A2 => gl_rom_n_637, A3 => gl_rom_n_633, A4 => gl_rom_n_630, ZN => gl_rom_n_1213);
  gl_rom_g35205 : ND4D0BWP7T port map(A1 => gl_rom_n_619, A2 => gl_rom_n_624, A3 => gl_rom_n_632, A4 => gl_rom_n_616, ZN => gl_rom_n_1212);
  gl_rom_g35206 : ND4D0BWP7T port map(A1 => gl_rom_n_625, A2 => gl_rom_n_631, A3 => gl_rom_n_629, A4 => gl_rom_n_626, ZN => gl_rom_n_1211);
  gl_rom_g35207 : ND4D0BWP7T port map(A1 => gl_rom_n_617, A2 => gl_rom_n_620, A3 => gl_rom_n_622, A4 => gl_rom_n_615, ZN => gl_rom_n_1210);
  gl_rom_g35208 : ND4D0BWP7T port map(A1 => gl_rom_n_609, A2 => gl_rom_n_621, A3 => gl_rom_n_618, A4 => gl_rom_n_614, ZN => gl_rom_n_1209);
  gl_rom_g35209 : ND4D0BWP7T port map(A1 => gl_rom_n_611, A2 => gl_rom_n_612, A3 => gl_rom_n_613, A4 => gl_rom_n_610, ZN => gl_rom_n_1208);
  gl_rom_g35210 : ND4D0BWP7T port map(A1 => gl_rom_n_596, A2 => gl_rom_n_581, A3 => gl_rom_n_600, A4 => gl_rom_n_588, ZN => gl_rom_n_1207);
  gl_rom_g35211 : ND4D0BWP7T port map(A1 => gl_rom_n_603, A2 => gl_rom_n_606, A3 => gl_rom_n_607, A4 => gl_rom_n_602, ZN => gl_rom_n_1206);
  gl_rom_g35212 : ND4D0BWP7T port map(A1 => gl_rom_n_605, A2 => gl_rom_n_598, A3 => gl_rom_n_601, A4 => gl_rom_n_593, ZN => gl_rom_n_1205);
  gl_rom_g35213 : ND4D0BWP7T port map(A1 => gl_rom_n_597, A2 => gl_rom_n_599, A3 => gl_rom_n_595, A4 => gl_rom_n_594, ZN => gl_rom_n_1204);
  gl_rom_g35214 : ND4D0BWP7T port map(A1 => gl_rom_n_585, A2 => gl_rom_n_579, A3 => gl_rom_n_591, A4 => gl_rom_n_584, ZN => gl_rom_n_1203);
  gl_rom_g35215 : ND4D0BWP7T port map(A1 => gl_rom_n_590, A2 => gl_rom_n_592, A3 => gl_rom_n_587, A4 => gl_rom_n_586, ZN => gl_rom_n_1202);
  gl_rom_g35216 : ND4D0BWP7T port map(A1 => gl_rom_n_582, A2 => gl_rom_n_583, A3 => gl_rom_n_580, A4 => gl_rom_n_578, ZN => gl_rom_n_1201);
  gl_rom_g35217 : ND4D0BWP7T port map(A1 => gl_rom_n_455, A2 => gl_rom_n_604, A3 => gl_rom_n_577, A4 => gl_rom_n_482, ZN => gl_rom_n_1200);
  gl_rom_g35218 : ND4D0BWP7T port map(A1 => gl_rom_n_514, A2 => gl_rom_n_545, A3 => gl_rom_n_575, A4 => gl_rom_n_490, ZN => gl_rom_n_1199);
  gl_rom_g35219 : ND4D0BWP7T port map(A1 => gl_rom_n_572, A2 => gl_rom_n_573, A3 => gl_rom_n_576, A4 => gl_rom_n_569, ZN => gl_rom_n_1198);
  gl_rom_g35220 : ND4D0BWP7T port map(A1 => gl_rom_n_568, A2 => gl_rom_n_542, A3 => gl_rom_n_558, A4 => gl_rom_n_529, ZN => gl_rom_n_1197);
  gl_rom_g35221 : ND4D0BWP7T port map(A1 => gl_rom_n_574, A2 => gl_rom_n_566, A3 => gl_rom_n_570, A4 => gl_rom_n_564, ZN => gl_rom_n_1196);
  gl_rom_g35222 : ND4D0BWP7T port map(A1 => gl_rom_n_554, A2 => gl_rom_n_561, A3 => gl_rom_n_571, A4 => gl_rom_n_551, ZN => gl_rom_n_1195);
  gl_rom_g35223 : ND4D0BWP7T port map(A1 => gl_rom_n_565, A2 => gl_rom_n_567, A3 => gl_rom_n_563, A4 => gl_rom_n_562, ZN => gl_rom_n_1194);
  gl_rom_g35224 : ND4D0BWP7T port map(A1 => gl_rom_n_556, A2 => gl_rom_n_548, A3 => gl_rom_n_560, A4 => gl_rom_n_552, ZN => gl_rom_n_1193);
  gl_rom_g35225 : ND4D0BWP7T port map(A1 => gl_rom_n_557, A2 => gl_rom_n_559, A3 => gl_rom_n_555, A4 => gl_rom_n_553, ZN => gl_rom_n_1192);
  gl_rom_g35226 : ND4D0BWP7T port map(A1 => gl_rom_n_911, A2 => gl_rom_n_756, A3 => gl_rom_n_862, A4 => gl_rom_n_641, ZN => gl_rom_n_1191);
  gl_rom_g35227 : ND4D0BWP7T port map(A1 => gl_rom_n_39, A2 => gl_rom_n_41, A3 => gl_rom_n_43, A4 => gl_rom_n_806, ZN => gl_rom_n_1190);
  gl_rom_g35228 : ND4D0BWP7T port map(A1 => gl_rom_n_543, A2 => gl_rom_n_544, A3 => gl_rom_n_539, A4 => gl_rom_n_537, ZN => gl_rom_n_1189);
  gl_rom_g35229 : ND4D0BWP7T port map(A1 => gl_rom_n_535, A2 => gl_rom_n_538, A3 => gl_rom_n_541, A4 => gl_rom_n_531, ZN => gl_rom_n_1188);
  gl_rom_g35230 : ND4D0BWP7T port map(A1 => gl_rom_n_534, A2 => gl_rom_n_530, A3 => gl_rom_n_536, A4 => gl_rom_n_532, ZN => gl_rom_n_1187);
  gl_rom_g35231 : ND4D0BWP7T port map(A1 => gl_rom_n_528, A2 => gl_rom_n_523, A3 => gl_rom_n_526, A4 => gl_rom_n_522, ZN => gl_rom_n_1186);
  gl_rom_g35232 : ND4D0BWP7T port map(A1 => gl_rom_n_517, A2 => gl_rom_n_525, A3 => gl_rom_n_524, A4 => gl_rom_n_519, ZN => gl_rom_n_1185);
  gl_rom_g35233 : ND4D0BWP7T port map(A1 => gl_rom_n_521, A2 => gl_rom_n_516, A3 => gl_rom_n_518, A4 => gl_rom_n_515, ZN => gl_rom_n_1184);
  gl_rom_g35234 : ND4D0BWP7T port map(A1 => gl_rom_n_498, A2 => gl_rom_n_476, A3 => gl_rom_n_510, A4 => gl_rom_n_480, ZN => gl_rom_n_1183);
  gl_rom_g35235 : ND4D0BWP7T port map(A1 => gl_rom_n_509, A2 => gl_rom_n_512, A3 => gl_rom_n_513, A4 => gl_rom_n_508, ZN => gl_rom_n_1182);
  gl_rom_g35236 : ND4D0BWP7T port map(A1 => gl_rom_n_511, A2 => gl_rom_n_504, A3 => gl_rom_n_507, A4 => gl_rom_n_501, ZN => gl_rom_n_1181);
  gl_rom_g35237 : ND4D0BWP7T port map(A1 => gl_rom_n_487, A2 => gl_rom_n_505, A3 => gl_rom_n_502, A4 => gl_rom_n_493, ZN => gl_rom_n_1180);
  gl_rom_g35238 : ND4D0BWP7T port map(A1 => gl_rom_n_500, A2 => gl_rom_n_503, A3 => gl_rom_n_506, A4 => gl_rom_n_499, ZN => gl_rom_n_1179);
  gl_rom_g35239 : ND4D0BWP7T port map(A1 => gl_rom_n_425, A2 => gl_rom_n_271, A3 => gl_rom_n_326, A4 => gl_rom_n_203, ZN => gl_rom_n_1178);
  gl_rom_g35240 : ND4D0BWP7T port map(A1 => gl_rom_n_488, A2 => gl_rom_n_492, A3 => gl_rom_n_496, A4 => gl_rom_n_485, ZN => gl_rom_n_1177);
  gl_rom_g35241 : ND4D0BWP7T port map(A1 => gl_rom_n_495, A2 => gl_rom_n_497, A3 => gl_rom_n_494, A4 => gl_rom_n_491, ZN => gl_rom_n_1176);
  gl_rom_g35242 : ND4D0BWP7T port map(A1 => gl_rom_n_484, A2 => gl_rom_n_486, A3 => gl_rom_n_489, A4 => gl_rom_n_483, ZN => gl_rom_n_1175);
  gl_rom_g35243 : ND4D0BWP7T port map(A1 => gl_rom_n_477, A2 => gl_rom_n_479, A3 => gl_rom_n_481, A4 => gl_rom_n_474, ZN => gl_rom_n_1174);
  gl_rom_g35244 : ND4D0BWP7T port map(A1 => gl_rom_n_478, A2 => gl_rom_n_469, A3 => gl_rom_n_475, A4 => gl_rom_n_467, ZN => gl_rom_n_1173);
  gl_rom_g35245 : ND4D0BWP7T port map(A1 => gl_rom_n_462, A2 => gl_rom_n_471, A3 => gl_rom_n_473, A4 => gl_rom_n_454, ZN => gl_rom_n_1172);
  gl_rom_g35246 : ND4D0BWP7T port map(A1 => gl_rom_n_466, A2 => gl_rom_n_472, A3 => gl_rom_n_470, A4 => gl_rom_n_468, ZN => gl_rom_n_1171);
  gl_rom_g35247 : ND4D0BWP7T port map(A1 => gl_rom_n_419, A2 => gl_rom_n_363, A3 => gl_rom_n_450, A4 => gl_rom_n_386, ZN => gl_rom_n_1170);
  gl_rom_g35248 : ND4D0BWP7T port map(A1 => gl_rom_n_464, A2 => gl_rom_n_457, A3 => gl_rom_n_460, A4 => gl_rom_n_452, ZN => gl_rom_n_1169);
  gl_rom_g35249 : ND4D0BWP7T port map(A1 => gl_rom_n_463, A2 => gl_rom_n_459, A3 => gl_rom_n_465, A4 => gl_rom_n_461, ZN => gl_rom_n_1168);
  gl_rom_g35250 : ND4D0BWP7T port map(A1 => gl_rom_n_458, A2 => gl_rom_n_453, A3 => gl_rom_n_456, A4 => gl_rom_n_451, ZN => gl_rom_n_1167);
  gl_rom_g35251 : ND4D0BWP7T port map(A1 => gl_rom_n_443, A2 => gl_rom_n_449, A3 => gl_rom_n_447, A4 => gl_rom_n_446, ZN => gl_rom_n_1166);
  gl_rom_g35252 : ND4D0BWP7T port map(A1 => gl_rom_n_401, A2 => gl_rom_n_445, A3 => gl_rom_n_432, A4 => gl_rom_n_416, ZN => gl_rom_n_1165);
  gl_rom_g35253 : ND4D0BWP7T port map(A1 => gl_rom_n_448, A2 => gl_rom_n_440, A3 => gl_rom_n_444, A4 => gl_rom_n_438, ZN => gl_rom_n_1164);
  gl_rom_g35254 : ND4D0BWP7T port map(A1 => gl_rom_n_435, A2 => gl_rom_n_424, A3 => gl_rom_n_442, A4 => gl_rom_n_428, ZN => gl_rom_n_1163);
  gl_rom_g35255 : ND4D0BWP7T port map(A1 => gl_rom_n_437, A2 => gl_rom_n_439, A3 => gl_rom_n_441, A4 => gl_rom_n_436, ZN => gl_rom_n_1162);
  gl_rom_g35256 : ND4D0BWP7T port map(A1 => gl_rom_n_430, A2 => gl_rom_n_434, A3 => gl_rom_n_426, A4 => gl_rom_n_421, ZN => gl_rom_n_1161);
  gl_rom_g35257 : ND4D0BWP7T port map(A1 => gl_rom_n_429, A2 => gl_rom_n_431, A3 => gl_rom_n_433, A4 => gl_rom_n_427, ZN => gl_rom_n_1160);
  gl_rom_g35258 : ND4D0BWP7T port map(A1 => gl_rom_n_420, A2 => gl_rom_n_422, A3 => gl_rom_n_423, A4 => gl_rom_n_418, ZN => gl_rom_n_1159);
  gl_rom_g35259 : ND4D0BWP7T port map(A1 => gl_rom_n_413, A2 => gl_rom_n_415, A3 => gl_rom_n_417, A4 => gl_rom_n_411, ZN => gl_rom_n_1158);
  gl_rom_g35260 : ND4D0BWP7T port map(A1 => gl_rom_n_410, A2 => gl_rom_n_414, A3 => gl_rom_n_407, A4 => gl_rom_n_406, ZN => gl_rom_n_1157);
  gl_rom_g35261 : ND4D0BWP7T port map(A1 => gl_rom_n_398, A2 => gl_rom_n_403, A3 => gl_rom_n_412, A4 => gl_rom_n_393, ZN => gl_rom_n_1156);
  gl_rom_g35262 : ND4D0BWP7T port map(A1 => gl_rom_n_409, A2 => gl_rom_n_405, A3 => gl_rom_n_408, A4 => gl_rom_n_404, ZN => gl_rom_n_1155);
  gl_rom_g35263 : ND4D0BWP7T port map(A1 => gl_rom_n_397, A2 => gl_rom_n_399, A3 => gl_rom_n_402, A4 => gl_rom_n_395, ZN => gl_rom_n_1154);
  gl_rom_g35264 : ND4D0BWP7T port map(A1 => gl_rom_n_392, A2 => gl_rom_n_396, A3 => gl_rom_n_400, A4 => gl_rom_n_390, ZN => gl_rom_n_1153);
  gl_rom_g35265 : ND4D0BWP7T port map(A1 => gl_rom_n_394, A2 => gl_rom_n_389, A3 => gl_rom_n_391, A4 => gl_rom_n_388, ZN => gl_rom_n_1152);
  gl_rom_g35266 : ND4D0BWP7T port map(A1 => gl_rom_n_370, A2 => gl_rom_n_384, A3 => gl_rom_n_353, A4 => gl_rom_n_342, ZN => gl_rom_n_1151);
  gl_rom_g35267 : ND4D0BWP7T port map(A1 => gl_rom_n_381, A2 => gl_rom_n_383, A3 => gl_rom_n_385, A4 => gl_rom_n_379, ZN => gl_rom_n_1150);
  gl_rom_g35268 : ND4D0BWP7T port map(A1 => gl_rom_n_382, A2 => gl_rom_n_376, A3 => gl_rom_n_380, A4 => gl_rom_n_373, ZN => gl_rom_n_1149);
  gl_rom_g35269 : ND4D0BWP7T port map(A1 => gl_rom_n_378, A2 => gl_rom_n_362, A3 => gl_rom_n_374, A4 => gl_rom_n_359, ZN => gl_rom_n_1148);
  gl_rom_g35270 : ND4D0BWP7T port map(A1 => gl_rom_n_372, A2 => gl_rom_n_375, A3 => gl_rom_n_377, A4 => gl_rom_n_371, ZN => gl_rom_n_1147);
  gl_rom_g35271 : ND4D0BWP7T port map(A1 => gl_rom_n_357, A2 => gl_rom_n_368, A3 => gl_rom_n_365, A4 => gl_rom_n_361, ZN => gl_rom_n_1146);
  gl_rom_g35272 : ND4D0BWP7T port map(A1 => gl_rom_n_366, A2 => gl_rom_n_367, A3 => gl_rom_n_369, A4 => gl_rom_n_364, ZN => gl_rom_n_1145);
  gl_rom_g35273 : ND4D0BWP7T port map(A1 => gl_rom_n_356, A2 => gl_rom_n_358, A3 => gl_rom_n_360, A4 => gl_rom_n_355, ZN => gl_rom_n_1144);
  gl_rom_g35274 : ND4D0BWP7T port map(A1 => gl_rom_n_329, A2 => gl_rom_n_350, A3 => gl_rom_n_341, A4 => gl_rom_n_331, ZN => gl_rom_n_1143);
  gl_rom_g35275 : ND4D0BWP7T port map(A1 => gl_rom_n_349, A2 => gl_rom_n_351, A3 => gl_rom_n_354, A4 => gl_rom_n_347, ZN => gl_rom_n_1142);
  gl_rom_g35276 : ND4D0BWP7T port map(A1 => gl_rom_n_348, A2 => gl_rom_n_339, A3 => gl_rom_n_352, A4 => gl_rom_n_343, ZN => gl_rom_n_1141);
  gl_rom_g35277 : ND4D0BWP7T port map(A1 => gl_rom_n_338, A2 => gl_rom_n_346, A3 => gl_rom_n_344, A4 => gl_rom_n_340, ZN => gl_rom_n_1140);
  gl_rom_g35278 : ND4D0BWP7T port map(A1 => gl_rom_n_257, A2 => gl_rom_n_345, A3 => gl_rom_n_289, A4 => gl_rom_n_265, ZN => gl_rom_n_1139);
  gl_rom_g35279 : ND4D0BWP7T port map(A1 => gl_rom_n_336, A2 => gl_rom_n_328, A3 => gl_rom_n_334, A4 => gl_rom_n_325, ZN => gl_rom_n_1138);
  gl_rom_g35280 : ND4D0BWP7T port map(A1 => gl_rom_n_333, A2 => gl_rom_n_335, A3 => gl_rom_n_337, A4 => gl_rom_n_332, ZN => gl_rom_n_1137);
  gl_rom_g35281 : ND4D0BWP7T port map(A1 => gl_rom_n_327, A2 => gl_rom_n_330, A3 => gl_rom_n_324, A4 => gl_rom_n_323, ZN => gl_rom_n_1136);
  gl_rom_g35282 : ND4D0BWP7T port map(A1 => gl_rom_n_288, A2 => gl_rom_n_302, A3 => gl_rom_n_322, A4 => gl_rom_n_279, ZN => gl_rom_n_1135);
  gl_rom_g35283 : ND4D0BWP7T port map(A1 => gl_rom_n_315, A2 => gl_rom_n_321, A3 => gl_rom_n_319, A4 => gl_rom_n_318, ZN => gl_rom_n_1134);
  gl_rom_g35284 : ND4D0BWP7T port map(A1 => gl_rom_n_317, A2 => gl_rom_n_298, A3 => gl_rom_n_309, A4 => gl_rom_n_293, ZN => gl_rom_n_1133);
  gl_rom_g35285 : ND4D0BWP7T port map(A1 => gl_rom_n_312, A2 => gl_rom_n_316, A3 => gl_rom_n_320, A4 => gl_rom_n_308, ZN => gl_rom_n_1132);
  gl_rom_g35286 : ND4D0BWP7T port map(A1 => gl_rom_n_304, A2 => gl_rom_n_313, A3 => gl_rom_n_314, A4 => gl_rom_n_301, ZN => gl_rom_n_1131);
  gl_rom_g35287 : ND4D0BWP7T port map(A1 => gl_rom_n_310, A2 => gl_rom_n_311, A3 => gl_rom_n_307, A4 => gl_rom_n_306, ZN => gl_rom_n_1130);
  gl_rom_g35288 : ND4D0BWP7T port map(A1 => gl_rom_n_299, A2 => gl_rom_n_305, A3 => gl_rom_n_303, A4 => gl_rom_n_300, ZN => gl_rom_n_1129);
  gl_rom_g35289 : ND4D0BWP7T port map(A1 => gl_rom_n_286, A2 => gl_rom_n_297, A3 => gl_rom_n_296, A4 => gl_rom_n_291, ZN => gl_rom_n_1128);
  gl_rom_g35290 : ND4D0BWP7T port map(A1 => gl_rom_n_292, A2 => gl_rom_n_550, A3 => gl_rom_n_295, A4 => gl_rom_n_290, ZN => gl_rom_n_1127);
  gl_rom_g35291 : ND4D0BWP7T port map(A1 => gl_rom_n_284, A2 => gl_rom_n_285, A3 => gl_rom_n_287, A4 => gl_rom_n_283, ZN => gl_rom_n_1126);
  gl_rom_g35292 : ND4D0BWP7T port map(A1 => gl_rom_n_282, A2 => gl_rom_n_270, A3 => gl_rom_n_281, A4 => gl_rom_n_262, ZN => gl_rom_n_1125);
  gl_rom_g35293 : ND4D0BWP7T port map(A1 => gl_rom_n_276, A2 => gl_rom_n_278, A3 => gl_rom_n_280, A4 => gl_rom_n_274, ZN => gl_rom_n_1124);
  gl_rom_g35294 : ND4D0BWP7T port map(A1 => gl_rom_n_275, A2 => gl_rom_n_277, A3 => gl_rom_n_269, A4 => gl_rom_n_266, ZN => gl_rom_n_1123);
  gl_rom_g35295 : ND4D0BWP7T port map(A1 => gl_rom_n_268, A2 => gl_rom_n_272, A3 => gl_rom_n_273, A4 => gl_rom_n_267, ZN => gl_rom_n_1122);
  gl_rom_g35296 : ND4D0BWP7T port map(A1 => gl_rom_n_254, A2 => gl_rom_n_259, A3 => gl_rom_n_261, A4 => gl_rom_n_250, ZN => gl_rom_n_1121);
  gl_rom_g35297 : ND4D0BWP7T port map(A1 => gl_rom_n_260, A2 => gl_rom_n_263, A3 => gl_rom_n_264, A4 => gl_rom_n_258, ZN => gl_rom_n_1120);
  gl_rom_g35298 : ND4D0BWP7T port map(A1 => gl_rom_n_252, A2 => gl_rom_n_255, A3 => gl_rom_n_256, A4 => gl_rom_n_251, ZN => gl_rom_n_1119);
  gl_rom_g35299 : ND4D0BWP7T port map(A1 => gl_rom_n_218, A2 => gl_rom_n_253, A3 => gl_rom_n_249, A4 => gl_rom_n_223, ZN => gl_rom_n_1118);
  gl_rom_g35300 : ND4D0BWP7T port map(A1 => gl_rom_n_243, A2 => gl_rom_n_248, A3 => gl_rom_n_247, A4 => gl_rom_n_245, ZN => gl_rom_n_1117);
  gl_rom_g35301 : ND4D0BWP7T port map(A1 => gl_rom_n_239, A2 => gl_rom_n_242, A3 => gl_rom_n_246, A4 => gl_rom_n_237, ZN => gl_rom_n_1116);
  gl_rom_g35302 : ND4D0BWP7T port map(A1 => gl_rom_n_235, A2 => gl_rom_n_227, A3 => gl_rom_n_244, A4 => gl_rom_n_231, ZN => gl_rom_n_1115);
  gl_rom_g35303 : ND4D0BWP7T port map(A1 => gl_rom_n_236, A2 => gl_rom_n_241, A3 => gl_rom_n_240, A4 => gl_rom_n_238, ZN => gl_rom_n_1114);
  gl_rom_g35304 : ND4D0BWP7T port map(A1 => gl_rom_n_228, A2 => gl_rom_n_232, A3 => gl_rom_n_225, A4 => gl_rom_n_222, ZN => gl_rom_n_1113);
  gl_rom_g35305 : ND4D0BWP7T port map(A1 => gl_rom_n_229, A2 => gl_rom_n_234, A3 => gl_rom_n_233, A4 => gl_rom_n_230, ZN => gl_rom_n_1112);
  gl_rom_g35306 : ND4D0BWP7T port map(A1 => gl_rom_n_220, A2 => gl_rom_n_226, A3 => gl_rom_n_224, A4 => gl_rom_n_221, ZN => gl_rom_n_1111);
  gl_rom_g35307 : ND4D0BWP7T port map(A1 => gl_rom_n_217, A2 => gl_rom_n_219, A3 => gl_rom_n_214, A4 => gl_rom_n_213, ZN => gl_rom_n_1110);
  gl_rom_g35308 : ND4D0BWP7T port map(A1 => gl_rom_n_216, A2 => gl_rom_n_199, A3 => gl_rom_n_211, A4 => gl_rom_n_193, ZN => gl_rom_n_1109);
  gl_rom_g35309 : ND4D0BWP7T port map(A1 => gl_rom_n_195, A2 => gl_rom_n_144, A3 => gl_rom_n_180, A4 => gl_rom_n_116, ZN => gl_rom_n_1108);
  gl_rom_g35310 : ND4D0BWP7T port map(A1 => gl_rom_n_208, A2 => gl_rom_n_212, A3 => gl_rom_n_215, A4 => gl_rom_n_205, ZN => gl_rom_n_1107);
  gl_rom_g35311 : ND4D0BWP7T port map(A1 => gl_rom_n_207, A2 => gl_rom_n_209, A3 => gl_rom_n_210, A4 => gl_rom_n_206, ZN => gl_rom_n_1106);
  gl_rom_g35312 : ND4D0BWP7T port map(A1 => gl_rom_n_189, A2 => gl_rom_n_201, A3 => gl_rom_n_197, A4 => gl_rom_n_191, ZN => gl_rom_n_1105);
  gl_rom_g35313 : ND4D0BWP7T port map(A1 => gl_rom_n_204, A2 => gl_rom_n_198, A3 => gl_rom_n_200, A4 => gl_rom_n_196, ZN => gl_rom_n_1104);
  gl_rom_g35314 : ND4D0BWP7T port map(A1 => gl_rom_n_192, A2 => gl_rom_n_188, A3 => gl_rom_n_194, A4 => gl_rom_n_190, ZN => gl_rom_n_1103);
  gl_rom_g35315 : ND4D0BWP7T port map(A1 => gl_rom_n_184, A2 => gl_rom_n_186, A3 => gl_rom_n_187, A4 => gl_rom_n_181, ZN => gl_rom_n_1102);
  gl_rom_g35316 : ND4D0BWP7T port map(A1 => gl_rom_n_178, A2 => gl_rom_n_163, A3 => gl_rom_n_183, A4 => gl_rom_n_169, ZN => gl_rom_n_1101);
  gl_rom_g35317 : ND4D0BWP7T port map(A1 => gl_rom_n_176, A2 => gl_rom_n_182, A3 => gl_rom_n_185, A4 => gl_rom_n_172, ZN => gl_rom_n_1100);
  gl_rom_g35318 : ND4D0BWP7T port map(A1 => gl_rom_n_140, A2 => gl_rom_n_175, A3 => gl_rom_n_171, A4 => gl_rom_n_151, ZN => gl_rom_n_1099);
  gl_rom_g35319 : ND4D0BWP7T port map(A1 => gl_rom_n_173, A2 => gl_rom_n_179, A3 => gl_rom_n_177, A4 => gl_rom_n_174, ZN => gl_rom_n_1098);
  gl_rom_g35320 : ND4D0BWP7T port map(A1 => gl_rom_n_165, A2 => gl_rom_n_167, A3 => gl_rom_n_170, A4 => gl_rom_n_164, ZN => gl_rom_n_1097);
  gl_rom_g35321 : ND4D0BWP7T port map(A1 => gl_rom_n_162, A2 => gl_rom_n_166, A3 => gl_rom_n_168, A4 => gl_rom_n_159, ZN => gl_rom_n_1096);
  gl_rom_g35322 : ND4D0BWP7T port map(A1 => gl_rom_n_161, A2 => gl_rom_n_158, A3 => gl_rom_n_160, A4 => gl_rom_n_157, ZN => gl_rom_n_1095);
  gl_rom_g35323 : ND4D0BWP7T port map(A1 => gl_rom_n_154, A2 => gl_rom_n_139, A3 => gl_rom_n_148, A4 => gl_rom_n_132, ZN => gl_rom_n_1094);
  gl_rom_g35324 : ND4D0BWP7T port map(A1 => gl_rom_n_152, A2 => gl_rom_n_155, A3 => gl_rom_n_156, A4 => gl_rom_n_150, ZN => gl_rom_n_1093);
  gl_rom_g35325 : ND4D0BWP7T port map(A1 => gl_rom_n_145, A2 => gl_rom_n_149, A3 => gl_rom_n_153, A4 => gl_rom_n_141, ZN => gl_rom_n_1092);
  gl_rom_g35326 : ND4D0BWP7T port map(A1 => gl_rom_n_142, A2 => gl_rom_n_147, A3 => gl_rom_n_146, A4 => gl_rom_n_143, ZN => gl_rom_n_1091);
  gl_rom_g35327 : ND4D0BWP7T port map(A1 => gl_rom_n_127, A2 => gl_rom_n_136, A3 => gl_rom_n_134, A4 => gl_rom_n_130, ZN => gl_rom_n_1090);
  gl_rom_g35328 : ND4D0BWP7T port map(A1 => gl_rom_n_138, A2 => gl_rom_n_135, A3 => gl_rom_n_137, A4 => gl_rom_n_133, ZN => gl_rom_n_1089);
  gl_rom_g35329 : ND4D0BWP7T port map(A1 => gl_rom_n_131, A2 => gl_rom_n_128, A3 => gl_rom_n_129, A4 => gl_rom_n_126, ZN => gl_rom_n_1088);
  gl_rom_g35330 : ND4D0BWP7T port map(A1 => gl_rom_n_93, A2 => gl_rom_n_1028, A3 => gl_rom_n_72, A4 => gl_rom_n_973, ZN => gl_rom_n_1087);
  gl_rom_g35331 : ND4D0BWP7T port map(A1 => gl_rom_n_125, A2 => gl_rom_n_121, A3 => gl_rom_n_124, A4 => gl_rom_n_120, ZN => gl_rom_n_1086);
  gl_rom_g35332 : ND4D0BWP7T port map(A1 => gl_rom_n_78, A2 => gl_rom_n_387, A3 => gl_rom_n_772, A4 => gl_rom_n_202, ZN => gl_rom_n_1085);
  gl_rom_g35333 : ND4D0BWP7T port map(A1 => gl_rom_n_75, A2 => gl_rom_n_119, A3 => gl_rom_n_109, A4 => gl_rom_n_91, ZN => gl_rom_n_1084);
  gl_rom_g35334 : ND4D0BWP7T port map(A1 => gl_rom_n_101, A2 => gl_rom_n_122, A3 => gl_rom_n_114, A4 => gl_rom_n_107, ZN => gl_rom_n_1083);
  gl_rom_g35335 : ND4D0BWP7T port map(A1 => gl_rom_n_113, A2 => gl_rom_n_118, A3 => gl_rom_n_123, A4 => gl_rom_n_112, ZN => gl_rom_n_1082);
  gl_rom_g35336 : ND4D0BWP7T port map(A1 => gl_rom_n_115, A2 => gl_rom_n_110, A3 => gl_rom_n_117, A4 => gl_rom_n_111, ZN => gl_rom_n_1081);
  gl_rom_g35337 : ND4D0BWP7T port map(A1 => gl_rom_n_99, A2 => gl_rom_n_104, A3 => gl_rom_n_106, A4 => gl_rom_n_97, ZN => gl_rom_n_1080);
  gl_rom_g35338 : ND4D0BWP7T port map(A1 => gl_rom_n_105, A2 => gl_rom_n_108, A3 => gl_rom_n_103, A4 => gl_rom_n_102, ZN => gl_rom_n_1079);
  gl_rom_g35339 : ND4D0BWP7T port map(A1 => gl_rom_n_96, A2 => gl_rom_n_98, A3 => gl_rom_n_100, A4 => gl_rom_n_95, ZN => gl_rom_n_1078);
  gl_rom_g35340 : ND4D0BWP7T port map(A1 => gl_rom_n_88, A2 => gl_rom_n_92, A3 => gl_rom_n_94, A4 => gl_rom_n_87, ZN => gl_rom_n_1077);
  gl_rom_g35341 : ND4D0BWP7T port map(A1 => gl_rom_n_89, A2 => gl_rom_n_77, A3 => gl_rom_n_85, A4 => gl_rom_n_68, ZN => gl_rom_n_1076);
  gl_rom_g35342 : ND4D0BWP7T port map(A1 => gl_rom_n_82, A2 => gl_rom_n_86, A3 => gl_rom_n_90, A4 => gl_rom_n_79, ZN => gl_rom_n_1075);
  gl_rom_g35343 : ND4D0BWP7T port map(A1 => gl_rom_n_81, A2 => gl_rom_n_83, A3 => gl_rom_n_84, A4 => gl_rom_n_80, ZN => gl_rom_n_1074);
  gl_rom_g35344 : ND4D0BWP7T port map(A1 => gl_rom_n_65, A2 => gl_rom_n_70, A3 => gl_rom_n_74, A4 => gl_rom_n_63, ZN => gl_rom_n_1073);
  gl_rom_g35345 : ND4D0BWP7T port map(A1 => gl_rom_n_73, A2 => gl_rom_n_76, A3 => gl_rom_n_71, A4 => gl_rom_n_69, ZN => gl_rom_n_1072);
  gl_rom_g35346 : ND4D0BWP7T port map(A1 => gl_rom_n_64, A2 => gl_rom_n_66, A3 => gl_rom_n_67, A4 => gl_rom_n_62, ZN => gl_rom_n_1071);
  gl_rom_g35347 : ND4D0BWP7T port map(A1 => gl_rom_n_55, A2 => gl_rom_n_61, A3 => gl_rom_n_60, A4 => gl_rom_n_57, ZN => gl_rom_n_1070);
  gl_rom_g35348 : ND4D0BWP7T port map(A1 => gl_rom_n_58, A2 => gl_rom_n_44, A3 => gl_rom_n_53, A4 => gl_rom_n_1055, ZN => gl_rom_n_1069);
  gl_rom_g35349 : ND4D0BWP7T port map(A1 => gl_rom_n_52, A2 => gl_rom_n_56, A3 => gl_rom_n_59, A4 => gl_rom_n_49, ZN => gl_rom_n_1068);
  gl_rom_g35350 : ND4D0BWP7T port map(A1 => gl_rom_n_1053, A2 => gl_rom_n_45, A3 => gl_rom_n_50, A4 => gl_rom_n_1042, ZN => gl_rom_n_1067);
  gl_rom_g35351 : ND4D0BWP7T port map(A1 => gl_rom_n_48, A2 => gl_rom_n_51, A3 => gl_rom_n_54, A4 => gl_rom_n_47, ZN => gl_rom_n_1066);
  gl_rom_g35352 : ND4D0BWP7T port map(A1 => gl_rom_n_46, A2 => gl_rom_n_1021, A3 => gl_rom_n_1054, A4 => gl_rom_n_988, ZN => gl_rom_n_1065);
  gl_rom_g35353 : ND4D0BWP7T port map(A1 => gl_rom_n_1061, A2 => gl_rom_n_40, A3 => gl_rom_n_42, A4 => gl_rom_n_1058, ZN => gl_rom_n_1064);
  gl_rom_g35354 : ND4D0BWP7T port map(A1 => gl_rom_n_527, A2 => gl_rom_n_533, A3 => gl_rom_n_540, A4 => gl_rom_n_520, ZN => gl_rom_n_1063);
  gl_rom_g35355 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_776(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_779(0), ZN => gl_rom_n_1062);
  gl_rom_g35356 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_385(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_389(0), ZN => gl_rom_n_1061);
  gl_rom_g35357 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_977(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_981(1), ZN => gl_rom_n_1060);
  gl_rom_g35358 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_980(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_982(1), ZN => gl_rom_n_1059);
  gl_rom_g35359 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_384(0), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_387(0), ZN => gl_rom_n_1058);
  gl_rom_g35360 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_978(1), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_979(1), ZN => gl_rom_n_1057);
  gl_rom_g35361 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_976(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_983(1), ZN => gl_rom_n_1056);
  gl_rom_g35362 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_712(0), B1 => FE_OFN19_gl_rom_n_21, B2 => gl_rom_rom_713(0), ZN => gl_rom_n_1055);
  gl_rom_g35363 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_956(0), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_958(0), ZN => gl_rom_n_1054);
  gl_rom_g35364 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_882(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_887(0), ZN => gl_rom_n_1053);
  gl_rom_g35365 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_706(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_711(0), ZN => gl_rom_n_1052);
  gl_rom_g35366 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_985(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_989(1), ZN => gl_rom_n_1051);
  gl_rom_g35367 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_988(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_990(1), ZN => gl_rom_n_1050);
  gl_rom_g35368 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_378(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_383(0), ZN => gl_rom_n_1049);
  gl_rom_g35369 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_986(1), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_987(1), ZN => gl_rom_n_1048);
  gl_rom_g35370 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_984(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_991(1), ZN => gl_rom_n_1047);
  gl_rom_g35371 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_708(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_710(0), ZN => gl_rom_n_1046);
  gl_rom_g35372 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_380(0), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_382(0), ZN => gl_rom_n_1045);
  gl_rom_g35373 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_994(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_999(1), ZN => gl_rom_n_1044);
  gl_rom_g35374 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_21, A2 => gl_rom_rom_993(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_997(1), ZN => gl_rom_n_1043);
  gl_rom_g35375 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_880(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_883(0), ZN => gl_rom_n_1042);
  gl_rom_g35376 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_22, A2 => gl_rom_rom_381(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_379(0), ZN => gl_rom_n_1041);
  gl_rom_g35377 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_996(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_998(1), ZN => gl_rom_n_1040);
  gl_rom_g35378 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_376(0), B1 => FE_OFN20_gl_rom_n_21, B2 => gl_rom_rom_377(0), ZN => gl_rom_n_1039);
  gl_rom_g35379 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_992(1), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_995(1), ZN => gl_rom_n_1038);
  gl_rom_g35380 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_1020(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_1023(1), ZN => gl_rom_n_1037);
  gl_rom_g35381 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_22, A2 => gl_rom_rom_709(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_707(0), ZN => gl_rom_n_1036);
  gl_rom_g35382 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_1018(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_1022(1), ZN => gl_rom_n_1035);
  gl_rom_g35383 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_362(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_367(0), ZN => gl_rom_n_1034);
  gl_rom_g35384 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_704(0), B1 => FE_OFN19_gl_rom_n_21, B2 => gl_rom_rom_705(0), ZN => gl_rom_n_1033);
  gl_rom_g35385 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_1017(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_1021(1), ZN => gl_rom_n_1032);
  gl_rom_g35386 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_1016(1), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_1019(1), ZN => gl_rom_n_1031);
  gl_rom_g35387 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_361(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_365(0), ZN => gl_rom_n_1030);
  gl_rom_g35388 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_1004(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_1007(1), ZN => gl_rom_n_1029);
  gl_rom_g35389 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_997(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_995(0), ZN => gl_rom_n_1028);
  gl_rom_g35390 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_1002(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_1006(1), ZN => gl_rom_n_1027);
  gl_rom_g35391 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_364(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_366(0), ZN => gl_rom_n_1026);
  gl_rom_g35392 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_360(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_363(0), ZN => gl_rom_n_1025);
  gl_rom_g35393 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_1001(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_1005(1), ZN => gl_rom_n_1024);
  gl_rom_g35394 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_1000(1), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_1003(1), ZN => gl_rom_n_1023);
  gl_rom_g35395 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_972(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_975(1), ZN => gl_rom_n_1022);
  gl_rom_g35396 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_22, A2 => gl_rom_rom_957(0), B1 => FE_OFN17_gl_rom_n_15, B2 => gl_rom_rom_955(0), ZN => gl_rom_n_1021);
  gl_rom_g35397 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_970(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_974(1), ZN => gl_rom_n_1020);
  gl_rom_g35398 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_370(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_375(0), ZN => gl_rom_n_1019);
  gl_rom_g35399 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_969(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_973(1), ZN => gl_rom_n_1018);
  gl_rom_g35400 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_852(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_855(0), ZN => gl_rom_n_1017);
  gl_rom_g35401 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_968(1), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_971(1), ZN => gl_rom_n_1016);
  gl_rom_g35402 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_372(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_374(0), ZN => gl_rom_n_1015);
  gl_rom_g35403 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_794(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_799(0), ZN => gl_rom_n_1014);
  gl_rom_g35404 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_964(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_967(1), ZN => gl_rom_n_1013);
  gl_rom_g35405 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_22, A2 => gl_rom_rom_373(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_371(0), ZN => gl_rom_n_1012);
  gl_rom_g35406 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_962(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_966(1), ZN => gl_rom_n_1011);
  gl_rom_g35407 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_850(0), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_854(0), ZN => gl_rom_n_1010);
  gl_rom_g35408 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_961(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_965(1), ZN => gl_rom_n_1009);
  gl_rom_g35409 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_960(1), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_963(1), ZN => gl_rom_n_1008);
  gl_rom_g35410 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_368(0), B1 => FE_OFN19_gl_rom_n_21, B2 => gl_rom_rom_369(0), ZN => gl_rom_n_1007);
  gl_rom_g35411 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_953(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_957(1), ZN => gl_rom_n_1006);
  gl_rom_g35412 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_21, A2 => gl_rom_rom_793(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_797(0), ZN => gl_rom_n_1005);
  gl_rom_g35413 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_796(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_798(0), ZN => gl_rom_n_1004);
  gl_rom_g35414 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_956(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_958(1), ZN => gl_rom_n_1003);
  gl_rom_g35415 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_338(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_343(0), ZN => gl_rom_n_1002);
  gl_rom_g35416 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_954(1), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_955(1), ZN => gl_rom_n_1001);
  gl_rom_g35417 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_340(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_342(0), ZN => gl_rom_n_1000);
  gl_rom_g35418 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_952(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_959(1), ZN => gl_rom_n_999);
  gl_rom_g35419 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_792(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_795(0), ZN => gl_rom_n_998);
  gl_rom_g35420 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_937(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_941(1), ZN => gl_rom_n_997);
  gl_rom_g35421 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_22, A2 => gl_rom_rom_341(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_339(0), ZN => gl_rom_n_996);
  gl_rom_g35422 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_940(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_942(1), ZN => gl_rom_n_995);
  gl_rom_g35423 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_938(1), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_939(1), ZN => gl_rom_n_994);
  gl_rom_g35424 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_336(0), B1 => FE_OFN19_gl_rom_n_21, B2 => gl_rom_rom_337(0), ZN => gl_rom_n_993);
  gl_rom_g35425 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_936(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_943(1), ZN => gl_rom_n_992);
  gl_rom_g35426 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_924(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_927(1), ZN => gl_rom_n_991);
  gl_rom_g35427 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_21, A2 => gl_rom_rom_849(0), B1 => FE_OFN11_gl_rom_n_22, B2 => gl_rom_rom_853(0), ZN => gl_rom_n_990);
  gl_rom_g35428 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_922(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_926(1), ZN => gl_rom_n_989);
  gl_rom_g35429 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_952(0), B1 => FE_OFN20_gl_rom_n_21, B2 => gl_rom_rom_953(0), ZN => gl_rom_n_988);
  gl_rom_g35430 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_346(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_351(0), ZN => gl_rom_n_987);
  gl_rom_g35431 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_921(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_925(1), ZN => gl_rom_n_986);
  gl_rom_g35432 : AOI22D0BWP7T port map(A1 => FE_OFN3_gl_rom_n_16, A2 => gl_rom_rom_806(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_805(0), ZN => gl_rom_n_985);
  gl_rom_g35433 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_920(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_923(1), ZN => gl_rom_n_984);
  gl_rom_g35434 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_348(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_350(0), ZN => gl_rom_n_983);
  gl_rom_g35435 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_848(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_851(0), ZN => gl_rom_n_982);
  gl_rom_g35436 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_930(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_935(1), ZN => gl_rom_n_981);
  gl_rom_g35437 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_929(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_933(1), ZN => gl_rom_n_980);
  gl_rom_g35438 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_22, A2 => gl_rom_rom_349(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_347(0), ZN => gl_rom_n_979);
  gl_rom_g35439 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_932(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_934(1), ZN => gl_rom_n_978);
  gl_rom_g35440 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_344(0), B1 => FE_OFN19_gl_rom_n_21, B2 => gl_rom_rom_345(0), ZN => gl_rom_n_977);
  gl_rom_g35441 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_928(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_931(1), ZN => gl_rom_n_976);
  gl_rom_g35442 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_804(0), B1 => FE_OFN19_gl_rom_n_21, B2 => gl_rom_rom_801(0), ZN => gl_rom_n_975);
  gl_rom_g35443 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_945(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_949(1), ZN => gl_rom_n_974);
  gl_rom_g35444 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_992(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_993(0), ZN => gl_rom_n_973);
  gl_rom_g35445 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_948(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_950(1), ZN => gl_rom_n_972);
  gl_rom_g35446 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_354(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_359(0), ZN => gl_rom_n_971);
  gl_rom_g35447 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_802(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_807(0), ZN => gl_rom_n_970);
  gl_rom_g35448 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_946(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_947(1), ZN => gl_rom_n_969);
  gl_rom_g35449 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_356(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_358(0), ZN => gl_rom_n_968);
  gl_rom_g35450 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_944(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_951(1), ZN => gl_rom_n_967);
  gl_rom_g35451 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_914(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_919(1), ZN => gl_rom_n_966);
  gl_rom_g35452 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_800(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_803(0), ZN => gl_rom_n_965);
  gl_rom_g35453 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_22, A2 => gl_rom_rom_357(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_355(0), ZN => gl_rom_n_964);
  gl_rom_g35454 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_913(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_917(1), ZN => gl_rom_n_963);
  gl_rom_g35455 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_352(0), B1 => FE_OFN19_gl_rom_n_21, B2 => gl_rom_rom_353(0), ZN => gl_rom_n_962);
  gl_rom_g35456 : AOI22D0BWP7T port map(A1 => FE_OFN0_gl_rom_n_16, A2 => gl_rom_rom_918(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_915(1), ZN => gl_rom_n_961);
  gl_rom_g35457 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_912(1), B1 => gl_rom_n_18, B2 => gl_rom_rom_916(1), ZN => gl_rom_n_960);
  gl_rom_g35458 : AOI22D0BWP7T port map(A1 => FE_OFN0_gl_rom_n_16, A2 => gl_rom_rom_910(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_909(1), ZN => gl_rom_n_959);
  gl_rom_g35459 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_908(1), B1 => FE_OFN22_gl_rom_n_21, B2 => gl_rom_rom_905(1), ZN => gl_rom_n_958);
  gl_rom_g35460 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_21, A2 => gl_rom_rom_329(0), B1 => FE_OFN11_gl_rom_n_22, B2 => gl_rom_rom_333(0), ZN => gl_rom_n_957);
  gl_rom_g35461 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_906(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_911(1), ZN => gl_rom_n_956);
  gl_rom_g35462 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_904(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_907(1), ZN => gl_rom_n_955);
  gl_rom_g35463 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_332(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_334(0), ZN => gl_rom_n_954);
  gl_rom_g35464 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_21, A2 => gl_rom_rom_817(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_821(0), ZN => gl_rom_n_953);
  gl_rom_g35465 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_938(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_943(0), ZN => gl_rom_n_952);
  gl_rom_g35466 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_898(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_903(1), ZN => gl_rom_n_951);
  gl_rom_g35467 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_890(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_895(0), ZN => gl_rom_n_950);
  gl_rom_g35468 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_330(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_331(0), ZN => gl_rom_n_949);
  gl_rom_g35469 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_897(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_901(1), ZN => gl_rom_n_948);
  gl_rom_g35470 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_820(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_822(0), ZN => gl_rom_n_947);
  gl_rom_g35471 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_328(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_335(0), ZN => gl_rom_n_946);
  gl_rom_g35472 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_900(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_902(1), ZN => gl_rom_n_945);
  gl_rom_g35473 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_896(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_899(1), ZN => gl_rom_n_944);
  gl_rom_g35474 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_892(0), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_894(0), ZN => gl_rom_n_943);
  gl_rom_g35475 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_700(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_703(1), ZN => gl_rom_n_942);
  gl_rom_g35476 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_322(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_327(0), ZN => gl_rom_n_941);
  gl_rom_g35477 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_698(1), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_702(1), ZN => gl_rom_n_940);
  gl_rom_g35478 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_818(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_819(0), ZN => gl_rom_n_939);
  gl_rom_g35479 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_697(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_701(1), ZN => gl_rom_n_938);
  gl_rom_g35480 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_696(1), B1 => FE_OFN17_gl_rom_n_15, B2 => gl_rom_rom_699(1), ZN => gl_rom_n_937);
  gl_rom_g35481 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_324(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_326(0), ZN => gl_rom_n_936);
  gl_rom_g35482 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_22, A2 => gl_rom_rom_325(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_323(0), ZN => gl_rom_n_935);
  gl_rom_g35483 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_684(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_687(1), ZN => gl_rom_n_934);
  gl_rom_g35484 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_816(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_823(0), ZN => gl_rom_n_933);
  gl_rom_g35485 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_682(1), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_686(1), ZN => gl_rom_n_932);
  gl_rom_g35486 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_320(0), B1 => FE_OFN19_gl_rom_n_21, B2 => gl_rom_rom_321(0), ZN => gl_rom_n_931);
  gl_rom_g35487 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_681(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_685(1), ZN => gl_rom_n_930);
  gl_rom_g35488 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_680(1), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_683(1), ZN => gl_rom_n_929);
  gl_rom_g35489 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_22, A2 => gl_rom_rom_893(0), B1 => FE_OFN17_gl_rom_n_15, B2 => gl_rom_rom_891(0), ZN => gl_rom_n_928);
  gl_rom_g35490 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_690(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_695(1), ZN => gl_rom_n_927);
  gl_rom_g35491 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_692(1), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_694(1), ZN => gl_rom_n_926);
  gl_rom_g35492 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_940(0), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_942(0), ZN => gl_rom_n_925);
  gl_rom_g35493 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_124(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_127(0), ZN => gl_rom_n_924);
  gl_rom_g35494 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_22, A2 => gl_rom_rom_693(1), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_691(1), ZN => gl_rom_n_923);
  gl_rom_g35495 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_688(1), B1 => FE_OFN22_gl_rom_n_21, B2 => gl_rom_rom_689(1), ZN => gl_rom_n_922);
  gl_rom_g35496 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_122(0), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_126(0), ZN => gl_rom_n_921);
  gl_rom_g35497 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_660(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_663(1), ZN => gl_rom_n_920);
  gl_rom_g35498 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_786(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_791(0), ZN => gl_rom_n_919);
  gl_rom_g35499 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_658(1), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_662(1), ZN => gl_rom_n_918);
  gl_rom_g35500 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_21, A2 => gl_rom_rom_785(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_789(0), ZN => gl_rom_n_917);
  gl_rom_g35501 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_121(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_125(0), ZN => gl_rom_n_916);
  gl_rom_g35502 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_120(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_123(0), ZN => gl_rom_n_915);
  gl_rom_g35503 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_657(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_661(1), ZN => gl_rom_n_914);
  gl_rom_g35504 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_656(1), B1 => FE_OFN17_gl_rom_n_15, B2 => gl_rom_rom_659(1), ZN => gl_rom_n_913);
  gl_rom_g35505 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_666(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_671(1), ZN => gl_rom_n_912);
  gl_rom_g35506 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_978(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_983(0), ZN => gl_rom_n_911);
  gl_rom_g35507 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_888(0), B1 => FE_OFN20_gl_rom_n_21, B2 => gl_rom_rom_889(0), ZN => gl_rom_n_910);
  gl_rom_g35508 : AOI22D0BWP7T port map(A1 => FE_OFN3_gl_rom_n_16, A2 => gl_rom_rom_790(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_787(0), ZN => gl_rom_n_909);
  gl_rom_g35509 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_665(1), B1 => FE_OFN11_gl_rom_n_22, B2 => gl_rom_rom_669(1), ZN => gl_rom_n_908);
  gl_rom_g35510 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_106(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_111(0), ZN => gl_rom_n_907);
  gl_rom_g35511 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_105(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_109(0), ZN => gl_rom_n_906);
  gl_rom_g35512 : AOI22D0BWP7T port map(A1 => FE_OFN1_gl_rom_n_16, A2 => gl_rom_rom_670(1), B1 => FE_OFN17_gl_rom_n_15, B2 => gl_rom_rom_667(1), ZN => gl_rom_n_905);
  gl_rom_g35513 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_664(1), B1 => FE_OFN5_gl_rom_n_18, B2 => gl_rom_rom_668(1), ZN => gl_rom_n_904);
  gl_rom_g35514 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_676(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_679(1), ZN => gl_rom_n_903);
  gl_rom_g35515 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_22, A2 => gl_rom_rom_941(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_939(0), ZN => gl_rom_n_902);
  gl_rom_g35516 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_784(0), B1 => FE_OFN6_gl_rom_n_18, B2 => gl_rom_rom_788(0), ZN => gl_rom_n_901);
  gl_rom_g35517 : AOI22D0BWP7T port map(A1 => FE_OFN1_gl_rom_n_16, A2 => gl_rom_rom_110(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_107(0), ZN => gl_rom_n_900);
  gl_rom_g35518 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_674(1), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_678(1), ZN => gl_rom_n_899);
  gl_rom_g35519 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_104(0), B1 => FE_OFN5_gl_rom_n_18, B2 => gl_rom_rom_108(0), ZN => gl_rom_n_898);
  gl_rom_g35520 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_673(1), B1 => FE_OFN11_gl_rom_n_22, B2 => gl_rom_rom_677(1), ZN => gl_rom_n_897);
  gl_rom_g35521 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_672(1), B1 => FE_OFN17_gl_rom_n_15, B2 => gl_rom_rom_675(1), ZN => gl_rom_n_896);
  gl_rom_g35522 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_652(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_655(1), ZN => gl_rom_n_895);
  gl_rom_g35523 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_650(1), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_654(1), ZN => gl_rom_n_894);
  gl_rom_g35524 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_874(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_879(0), ZN => gl_rom_n_893);
  gl_rom_g35525 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_114(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_119(0), ZN => gl_rom_n_892);
  gl_rom_g35526 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_649(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_653(1), ZN => gl_rom_n_891);
  gl_rom_g35527 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_116(0), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_118(0), ZN => gl_rom_n_890);
  gl_rom_g35528 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_648(1), B1 => FE_OFN17_gl_rom_n_15, B2 => gl_rom_rom_651(1), ZN => gl_rom_n_889);
  gl_rom_g35529 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_21, A2 => gl_rom_rom_825(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_829(0), ZN => gl_rom_n_888);
  gl_rom_g35530 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_828(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_830(0), ZN => gl_rom_n_887);
  gl_rom_g35531 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_642(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_647(1), ZN => gl_rom_n_886);
  gl_rom_g35532 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_22, A2 => gl_rom_rom_117(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_115(0), ZN => gl_rom_n_885);
  gl_rom_g35533 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_641(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_645(1), ZN => gl_rom_n_884);
  gl_rom_g35534 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_644(1), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_646(1), ZN => gl_rom_n_883);
  gl_rom_g35535 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_640(1), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_643(1), ZN => gl_rom_n_882);
  gl_rom_g35536 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_569(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_573(1), ZN => gl_rom_n_881);
  gl_rom_g35537 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_112(0), B1 => FE_OFN20_gl_rom_n_21, B2 => gl_rom_rom_113(0), ZN => gl_rom_n_880);
  gl_rom_g35538 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_873(0), B1 => FE_OFN11_gl_rom_n_22, B2 => gl_rom_rom_877(0), ZN => gl_rom_n_879);
  gl_rom_g35539 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_82(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_87(0), ZN => gl_rom_n_878);
  gl_rom_g35540 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_572(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_574(1), ZN => gl_rom_n_877);
  gl_rom_g35541 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_826(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_827(0), ZN => gl_rom_n_876);
  gl_rom_g35542 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_570(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_571(1), ZN => gl_rom_n_875);
  gl_rom_g35543 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_84(0), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_86(0), ZN => gl_rom_n_874);
  gl_rom_g35544 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_568(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_575(1), ZN => gl_rom_n_873);
  gl_rom_g35545 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_824(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_831(0), ZN => gl_rom_n_872);
  gl_rom_g35546 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_22, A2 => gl_rom_rom_85(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_83(0), ZN => gl_rom_n_871);
  gl_rom_g35547 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_554(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_559(1), ZN => gl_rom_n_870);
  gl_rom_g35548 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_21, A2 => gl_rom_rom_553(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_557(1), ZN => gl_rom_n_869);
  gl_rom_g35549 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_556(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_558(1), ZN => gl_rom_n_868);
  gl_rom_g35550 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_80(0), B1 => FE_OFN20_gl_rom_n_21, B2 => gl_rom_rom_81(0), ZN => gl_rom_n_867);
  gl_rom_g35551 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_552(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_555(1), ZN => gl_rom_n_866);
  gl_rom_g35552 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_936(0), B1 => FE_OFN20_gl_rom_n_21, B2 => gl_rom_rom_937(0), ZN => gl_rom_n_865);
  gl_rom_g35553 : AOI22D0BWP7T port map(A1 => FE_OFN1_gl_rom_n_16, A2 => gl_rom_rom_878(0), B1 => FE_OFN17_gl_rom_n_15, B2 => gl_rom_rom_875(0), ZN => gl_rom_n_864);
  gl_rom_g35554 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_564(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_567(1), ZN => gl_rom_n_863);
  gl_rom_g35555 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_980(0), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_982(0), ZN => gl_rom_n_862);
  gl_rom_g35556 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_1018(0), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_1023(0), ZN => gl_rom_n_861);
  gl_rom_g35557 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_562(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_566(1), ZN => gl_rom_n_860);
  gl_rom_g35558 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_90(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_95(0), ZN => gl_rom_n_859);
  gl_rom_g35559 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_810(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_815(0), ZN => gl_rom_n_858);
  gl_rom_g35560 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_21, A2 => gl_rom_rom_561(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_565(1), ZN => gl_rom_n_857);
  gl_rom_g35561 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_92(0), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_94(0), ZN => gl_rom_n_856);
  gl_rom_g35562 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_560(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_563(1), ZN => gl_rom_n_855);
  gl_rom_g35563 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_532(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_535(1), ZN => gl_rom_n_854);
  gl_rom_g35564 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_22, A2 => gl_rom_rom_93(0), B1 => FE_OFN17_gl_rom_n_15, B2 => gl_rom_rom_91(0), ZN => gl_rom_n_853);
  gl_rom_g35565 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_530(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_534(1), ZN => gl_rom_n_852);
  gl_rom_g35566 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_21, A2 => gl_rom_rom_809(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_813(0), ZN => gl_rom_n_851);
  gl_rom_g35567 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_21, A2 => gl_rom_rom_529(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_533(1), ZN => gl_rom_n_850);
  gl_rom_g35568 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_528(1), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_531(1), ZN => gl_rom_n_849);
  gl_rom_g35569 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_88(0), B1 => FE_OFN20_gl_rom_n_21, B2 => gl_rom_rom_89(0), ZN => gl_rom_n_848);
  gl_rom_g35570 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_540(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_543(1), ZN => gl_rom_n_847);
  gl_rom_g35571 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_872(0), B1 => FE_OFN5_gl_rom_n_18, B2 => gl_rom_rom_876(0), ZN => gl_rom_n_846);
  gl_rom_g35572 : AOI22D0BWP7T port map(A1 => FE_OFN3_gl_rom_n_16, A2 => gl_rom_rom_814(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_811(0), ZN => gl_rom_n_845);
  gl_rom_g35573 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_100(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_103(0), ZN => gl_rom_n_844);
  gl_rom_g35574 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_538(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_542(1), ZN => gl_rom_n_843);
  gl_rom_g35575 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_98(0), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_102(0), ZN => gl_rom_n_842);
  gl_rom_g35576 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_21, A2 => gl_rom_rom_537(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_541(1), ZN => gl_rom_n_841);
  gl_rom_g35577 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_536(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_539(1), ZN => gl_rom_n_840);
  gl_rom_g35578 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_548(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_551(1), ZN => gl_rom_n_839);
  gl_rom_g35579 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_808(0), B1 => FE_OFN6_gl_rom_n_18, B2 => gl_rom_rom_812(0), ZN => gl_rom_n_838);
  gl_rom_g35580 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_97(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_101(0), ZN => gl_rom_n_837);
  gl_rom_g35581 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_546(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_550(1), ZN => gl_rom_n_836);
  gl_rom_g35582 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_96(0), B1 => FE_OFN17_gl_rom_n_15, B2 => gl_rom_rom_99(0), ZN => gl_rom_n_835);
  gl_rom_g35583 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_21, A2 => gl_rom_rom_545(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_549(1), ZN => gl_rom_n_834);
  gl_rom_g35584 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_544(1), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_547(1), ZN => gl_rom_n_833);
  gl_rom_g35585 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_524(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_527(1), ZN => gl_rom_n_832);
  gl_rom_g35586 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_522(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_526(1), ZN => gl_rom_n_831);
  gl_rom_g35587 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_74(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_79(0), ZN => gl_rom_n_830);
  gl_rom_g35588 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_842(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_847(0), ZN => gl_rom_n_829);
  gl_rom_g35589 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_21, A2 => gl_rom_rom_521(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_525(1), ZN => gl_rom_n_828);
  gl_rom_g35590 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_778(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_783(0), ZN => gl_rom_n_827);
  gl_rom_g35591 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_520(1), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_523(1), ZN => gl_rom_n_826);
  gl_rom_g35592 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_73(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_77(0), ZN => gl_rom_n_825);
  gl_rom_g35593 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_946(0), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_951(0), ZN => gl_rom_n_824);
  gl_rom_g35594 : AOI22D0BWP7T port map(A1 => FE_OFN0_gl_rom_n_16, A2 => gl_rom_rom_518(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_517(1), ZN => gl_rom_n_823);
  gl_rom_g35595 : AOI22D0BWP7T port map(A1 => FE_OFN1_gl_rom_n_16, A2 => gl_rom_rom_78(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_75(0), ZN => gl_rom_n_822);
  gl_rom_g35596 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_516(1), B1 => FE_OFN23_gl_rom_n_21, B2 => gl_rom_rom_513(1), ZN => gl_rom_n_821);
  gl_rom_g35597 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_72(0), B1 => FE_OFN6_gl_rom_n_18, B2 => gl_rom_rom_76(0), ZN => gl_rom_n_820);
  gl_rom_g35598 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_514(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_519(1), ZN => gl_rom_n_819);
  gl_rom_g35599 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_512(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_515(1), ZN => gl_rom_n_818);
  gl_rom_g35600 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_21, A2 => gl_rom_rom_777(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_781(0), ZN => gl_rom_n_817);
  gl_rom_g35601 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_1017(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_1021(0), ZN => gl_rom_n_816);
  gl_rom_g35602 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_66(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_71(0), ZN => gl_rom_n_815);
  gl_rom_g35603 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_780(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_782(0), ZN => gl_rom_n_814);
  gl_rom_g35604 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_498(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_503(1), ZN => gl_rom_n_813);
  gl_rom_g35605 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_497(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_501(1), ZN => gl_rom_n_812);
  gl_rom_g35606 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_21, A2 => gl_rom_rom_841(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_845(0), ZN => gl_rom_n_811);
  gl_rom_g35607 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_68(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_70(0), ZN => gl_rom_n_810);
  gl_rom_g35608 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_500(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_502(1), ZN => gl_rom_n_809);
  gl_rom_g35609 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_496(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_499(1), ZN => gl_rom_n_808);
  gl_rom_g35610 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_22, A2 => gl_rom_rom_69(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_67(0), ZN => gl_rom_n_807);
  gl_rom_g35611 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_1008(1), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_1011(1), ZN => gl_rom_n_806);
  gl_rom_g35612 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_470(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_469(1), ZN => gl_rom_n_805);
  gl_rom_g35613 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_468(1), B1 => FE_OFN22_gl_rom_n_21, B2 => gl_rom_rom_465(1), ZN => gl_rom_n_804);
  gl_rom_g35614 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_64(0), B1 => FE_OFN20_gl_rom_n_21, B2 => gl_rom_rom_65(0), ZN => gl_rom_n_803);
  gl_rom_g35615 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_466(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_471(1), ZN => gl_rom_n_802);
  gl_rom_g35616 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_464(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_467(1), ZN => gl_rom_n_801);
  gl_rom_g35617 : AOI22D0BWP7T port map(A1 => FE_OFN1_gl_rom_n_16, A2 => gl_rom_rom_846(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_843(0), ZN => gl_rom_n_800);
  gl_rom_g35618 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_474(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_479(1), ZN => gl_rom_n_799);
  gl_rom_g35619 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_945(0), B1 => FE_OFN11_gl_rom_n_22, B2 => gl_rom_rom_949(0), ZN => gl_rom_n_798);
  gl_rom_g35620 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_770(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_775(0), ZN => gl_rom_n_797);
  gl_rom_g35621 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_476(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_478(1), ZN => gl_rom_n_796);
  gl_rom_g35622 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_21, A2 => gl_rom_rom_217(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_221(0), ZN => gl_rom_n_795);
  gl_rom_g35623 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_22, A2 => gl_rom_rom_477(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_475(1), ZN => gl_rom_n_794);
  gl_rom_g35624 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_472(1), B1 => FE_OFN22_gl_rom_n_21, B2 => gl_rom_rom_473(1), ZN => gl_rom_n_793);
  gl_rom_g35625 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_220(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_222(0), ZN => gl_rom_n_792);
  gl_rom_g35626 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_21, A2 => gl_rom_rom_769(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_773(0), ZN => gl_rom_n_791);
  gl_rom_g35627 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_484(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_487(1), ZN => gl_rom_n_790);
  gl_rom_g35628 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_482(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_486(1), ZN => gl_rom_n_789);
  gl_rom_g35629 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_218(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_219(0), ZN => gl_rom_n_788);
  gl_rom_g35630 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_481(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_485(1), ZN => gl_rom_n_787);
  gl_rom_g35631 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_480(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_483(1), ZN => gl_rom_n_786);
  gl_rom_g35632 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_216(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_223(0), ZN => gl_rom_n_785);
  gl_rom_g35633 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_506(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_511(1), ZN => gl_rom_n_784);
  gl_rom_g35634 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_840(0), B1 => FE_OFN6_gl_rom_n_18, B2 => gl_rom_rom_844(0), ZN => gl_rom_n_783);
  gl_rom_g35635 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_772(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_774(0), ZN => gl_rom_n_782);
  gl_rom_g35636 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_21, A2 => gl_rom_rom_225(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_229(0), ZN => gl_rom_n_781);
  gl_rom_g35637 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_508(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_510(1), ZN => gl_rom_n_780);
  gl_rom_g35638 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_768(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_771(0), ZN => gl_rom_n_779);
  gl_rom_g35639 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_22, A2 => gl_rom_rom_509(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_507(1), ZN => gl_rom_n_778);
  gl_rom_g35640 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_228(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_230(0), ZN => gl_rom_n_777);
  gl_rom_g35641 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_504(1), B1 => FE_OFN22_gl_rom_n_21, B2 => gl_rom_rom_505(1), ZN => gl_rom_n_776);
  gl_rom_g35642 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_494(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_493(1), ZN => gl_rom_n_775);
  gl_rom_g35643 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_226(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_227(0), ZN => gl_rom_n_774);
  gl_rom_g35644 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_492(1), B1 => FE_OFN22_gl_rom_n_21, B2 => gl_rom_rom_489(1), ZN => gl_rom_n_773);
  gl_rom_g35645 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_1012(0), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_1014(0), ZN => gl_rom_n_772);
  gl_rom_g35646 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_490(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_495(1), ZN => gl_rom_n_771);
  gl_rom_g35647 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_224(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_231(0), ZN => gl_rom_n_770);
  gl_rom_g35648 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_488(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_491(1), ZN => gl_rom_n_769);
  gl_rom_g35649 : AOI22D0BWP7T port map(A1 => FE_OFN0_gl_rom_n_16, A2 => gl_rom_rom_950(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_947(0), ZN => gl_rom_n_768);
  gl_rom_g35650 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_834(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_839(0), ZN => gl_rom_n_767);
  gl_rom_g35651 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_458(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_463(1), ZN => gl_rom_n_766);
  gl_rom_g35652 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_457(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_461(1), ZN => gl_rom_n_765);
  gl_rom_g35653 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_242(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_247(0), ZN => gl_rom_n_764);
  gl_rom_g35654 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_460(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_462(1), ZN => gl_rom_n_763);
  gl_rom_g35655 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_456(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_459(1), ZN => gl_rom_n_762);
  gl_rom_g35656 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_21, A2 => gl_rom_rom_241(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_245(0), ZN => gl_rom_n_761);
  gl_rom_g35657 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_700(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_703(0), ZN => gl_rom_n_760);
  gl_rom_g35658 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_454(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_453(1), ZN => gl_rom_n_759);
  gl_rom_g35659 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_244(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_246(0), ZN => gl_rom_n_758);
  gl_rom_g35660 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_452(1), B1 => FE_OFN22_gl_rom_n_21, B2 => gl_rom_rom_449(1), ZN => gl_rom_n_757);
  gl_rom_g35661 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_981(0), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_979(0), ZN => gl_rom_n_756);
  gl_rom_g35662 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_450(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_455(1), ZN => gl_rom_n_755);
  gl_rom_g35663 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_240(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_243(0), ZN => gl_rom_n_754);
  gl_rom_g35664 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_448(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_451(1), ZN => gl_rom_n_753);
  gl_rom_g35665 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_833(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_837(0), ZN => gl_rom_n_752);
  gl_rom_g35666 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_698(0), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_702(0), ZN => gl_rom_n_751);
  gl_rom_g35667 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_442(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_447(1), ZN => gl_rom_n_750);
  gl_rom_g35668 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_212(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_215(0), ZN => gl_rom_n_749);
  gl_rom_g35669 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_444(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_446(1), ZN => gl_rom_n_748);
  gl_rom_g35670 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_210(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_214(0), ZN => gl_rom_n_747);
  gl_rom_g35671 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_22, A2 => gl_rom_rom_445(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_443(1), ZN => gl_rom_n_746);
  gl_rom_g35672 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_440(1), B1 => FE_OFN22_gl_rom_n_21, B2 => gl_rom_rom_441(1), ZN => gl_rom_n_745);
  gl_rom_g35673 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_697(0), B1 => FE_OFN11_gl_rom_n_22, B2 => gl_rom_rom_701(0), ZN => gl_rom_n_744);
  gl_rom_g35674 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_1020(0), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_1022(0), ZN => gl_rom_n_743);
  gl_rom_g35675 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_944(0), B1 => FE_OFN7_gl_rom_n_18, B2 => gl_rom_rom_948(0), ZN => gl_rom_n_742);
  gl_rom_g35676 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_426(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_431(1), ZN => gl_rom_n_741);
  gl_rom_g35677 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_21, A2 => gl_rom_rom_209(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_213(0), ZN => gl_rom_n_740);
  gl_rom_g35678 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_425(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_429(1), ZN => gl_rom_n_739);
  gl_rom_g35679 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_428(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_430(1), ZN => gl_rom_n_738);
  gl_rom_g35680 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_424(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_427(1), ZN => gl_rom_n_737);
  gl_rom_g35681 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_208(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_211(0), ZN => gl_rom_n_736);
  gl_rom_g35682 : AOI22D0BWP7T port map(A1 => FE_OFN1_gl_rom_n_16, A2 => gl_rom_rom_838(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_835(0), ZN => gl_rom_n_735);
  gl_rom_g35683 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_410(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_415(1), ZN => gl_rom_n_734);
  gl_rom_g35684 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_409(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_413(1), ZN => gl_rom_n_733);
  gl_rom_g35685 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_696(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_699(0), ZN => gl_rom_n_732);
  gl_rom_g35686 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_252(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_255(0), ZN => gl_rom_n_731);
  gl_rom_g35687 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_412(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_414(1), ZN => gl_rom_n_730);
  gl_rom_g35688 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_250(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_254(0), ZN => gl_rom_n_729);
  gl_rom_g35689 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_408(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_411(1), ZN => gl_rom_n_728);
  gl_rom_g35690 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_681(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_685(0), ZN => gl_rom_n_727);
  gl_rom_g35691 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_832(0), B1 => FE_OFN6_gl_rom_n_18, B2 => gl_rom_rom_836(0), ZN => gl_rom_n_726);
  gl_rom_g35692 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_420(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_423(1), ZN => gl_rom_n_725);
  gl_rom_g35693 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_21, A2 => gl_rom_rom_249(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_253(0), ZN => gl_rom_n_724);
  gl_rom_g35694 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_418(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_422(1), ZN => gl_rom_n_723);
  gl_rom_g35695 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_684(0), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_686(0), ZN => gl_rom_n_722);
  gl_rom_g35696 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_417(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_421(1), ZN => gl_rom_n_721);
  gl_rom_g35697 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_416(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_419(1), ZN => gl_rom_n_720);
  gl_rom_g35698 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_248(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_251(0), ZN => gl_rom_n_719);
  gl_rom_g35699 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_438(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_437(1), ZN => gl_rom_n_718);
  gl_rom_g35700 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_436(1), B1 => FE_OFN22_gl_rom_n_21, B2 => gl_rom_rom_433(1), ZN => gl_rom_n_717);
  gl_rom_g35701 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_21, A2 => gl_rom_rom_233(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_237(0), ZN => gl_rom_n_716);
  gl_rom_g35702 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_434(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_439(1), ZN => gl_rom_n_715);
  gl_rom_g35703 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_236(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_238(0), ZN => gl_rom_n_714);
  gl_rom_g35704 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_432(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_435(1), ZN => gl_rom_n_713);
  gl_rom_g35705 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_682(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_683(0), ZN => gl_rom_n_712);
  gl_rom_g35706 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_402(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_407(1), ZN => gl_rom_n_711);
  gl_rom_g35707 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_234(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_235(0), ZN => gl_rom_n_710);
  gl_rom_g35708 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_401(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_405(1), ZN => gl_rom_n_709);
  gl_rom_g35709 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_680(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_687(0), ZN => gl_rom_n_708);
  gl_rom_g35710 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_404(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_406(1), ZN => gl_rom_n_707);
  gl_rom_g35711 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_1016(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_1019(0), ZN => gl_rom_n_706);
  gl_rom_g35712 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_232(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_239(0), ZN => gl_rom_n_705);
  gl_rom_g35713 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_400(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_403(1), ZN => gl_rom_n_704);
  gl_rom_g35714 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_914(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_919(0), ZN => gl_rom_n_703);
  gl_rom_g35715 : AOI22D0BWP7T port map(A1 => gl_rom_n_16, A2 => gl_rom_rom_398(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_397(1), ZN => gl_rom_n_702);
  gl_rom_g35716 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_396(1), B1 => FE_OFN22_gl_rom_n_21, B2 => gl_rom_rom_393(1), ZN => gl_rom_n_701);
  gl_rom_g35717 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_21, A2 => gl_rom_rom_201(0), B1 => FE_OFN11_gl_rom_n_22, B2 => gl_rom_rom_205(0), ZN => gl_rom_n_700);
  gl_rom_g35718 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_394(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_399(1), ZN => gl_rom_n_699);
  gl_rom_g35719 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_916(0), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_918(0), ZN => gl_rom_n_698);
  gl_rom_g35720 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_204(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_206(0), ZN => gl_rom_n_697);
  gl_rom_g35721 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_392(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_395(1), ZN => gl_rom_n_696);
  gl_rom_g35722 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_666(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_671(0), ZN => gl_rom_n_695);
  gl_rom_g35723 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_388(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_391(1), ZN => gl_rom_n_694);
  gl_rom_g35724 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_634(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_639(0), ZN => gl_rom_n_693);
  gl_rom_g35725 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_386(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_390(1), ZN => gl_rom_n_692);
  gl_rom_g35726 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_202(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_203(0), ZN => gl_rom_n_691);
  gl_rom_g35727 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_385(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_389(1), ZN => gl_rom_n_690);
  gl_rom_g35728 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_668(0), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_670(0), ZN => gl_rom_n_689);
  gl_rom_g35729 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_200(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_207(0), ZN => gl_rom_n_688);
  gl_rom_g35730 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_384(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_387(1), ZN => gl_rom_n_687);
  gl_rom_g35731 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_21, A2 => gl_rom_rom_193(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_197(0), ZN => gl_rom_n_686);
  gl_rom_g35732 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_249(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_253(1), ZN => gl_rom_n_685);
  gl_rom_g35733 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_252(1), B1 => FE_OFN4_gl_rom_n_16, B2 => gl_rom_rom_254(1), ZN => gl_rom_n_684);
  gl_rom_g35734 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_22, A2 => gl_rom_rom_669(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_667(0), ZN => gl_rom_n_683);
  gl_rom_g35735 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_196(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_198(0), ZN => gl_rom_n_682);
  gl_rom_g35736 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_250(1), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_251(1), ZN => gl_rom_n_681);
  gl_rom_g35737 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_248(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_255(1), ZN => gl_rom_n_680);
  gl_rom_g35738 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_636(0), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_638(0), ZN => gl_rom_n_679);
  gl_rom_g35739 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_194(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_195(0), ZN => gl_rom_n_678);
  gl_rom_g35740 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_234(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_239(1), ZN => gl_rom_n_677);
  gl_rom_g35741 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_233(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_237(1), ZN => gl_rom_n_676);
  gl_rom_g35742 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_192(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_199(0), ZN => gl_rom_n_675);
  gl_rom_g35743 : AOI22D0BWP7T port map(A1 => FE_OFN4_gl_rom_n_16, A2 => gl_rom_rom_238(1), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_235(1), ZN => gl_rom_n_674);
  gl_rom_g35744 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_232(1), B1 => FE_OFN7_gl_rom_n_18, B2 => gl_rom_rom_236(1), ZN => gl_rom_n_673);
  gl_rom_g35745 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_664(0), B1 => FE_OFN20_gl_rom_n_21, B2 => gl_rom_rom_665(0), ZN => gl_rom_n_672);
  gl_rom_g35746 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_241(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_245(1), ZN => gl_rom_n_671);
  gl_rom_g35747 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_244(1), B1 => FE_OFN4_gl_rom_n_16, B2 => gl_rom_rom_246(1), ZN => gl_rom_n_670);
  gl_rom_g35748 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_22, A2 => gl_rom_rom_637(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_635(0), ZN => gl_rom_n_669);
  gl_rom_g35749 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_316(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_319(0), ZN => gl_rom_n_668);
  gl_rom_g35750 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_242(1), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_243(1), ZN => gl_rom_n_667);
  gl_rom_g35751 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_240(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_247(1), ZN => gl_rom_n_666);
  gl_rom_g35752 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_674(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_679(0), ZN => gl_rom_n_665);
  gl_rom_g35753 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_314(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_318(0), ZN => gl_rom_n_664);
  gl_rom_g35754 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_676(0), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_678(0), ZN => gl_rom_n_663);
  gl_rom_g35755 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_212(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_215(1), ZN => gl_rom_n_662);
  gl_rom_g35756 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_210(1), B1 => FE_OFN4_gl_rom_n_16, B2 => gl_rom_rom_214(1), ZN => gl_rom_n_661);
  gl_rom_g35757 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_21, A2 => gl_rom_rom_313(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_317(0), ZN => gl_rom_n_660);
  gl_rom_g35758 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_209(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_213(1), ZN => gl_rom_n_659);
  gl_rom_g35759 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_208(1), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_211(1), ZN => gl_rom_n_658);
  gl_rom_g35760 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_312(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_315(0), ZN => gl_rom_n_657);
  gl_rom_g35761 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_218(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_223(1), ZN => gl_rom_n_656);
  gl_rom_g35762 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_22, A2 => gl_rom_rom_677(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_675(0), ZN => gl_rom_n_655);
  gl_rom_g35763 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_21, A2 => gl_rom_rom_217(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_221(1), ZN => gl_rom_n_654);
  gl_rom_g35764 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_300(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_303(0), ZN => gl_rom_n_653);
  gl_rom_g35765 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_632(0), B1 => FE_OFN20_gl_rom_n_21, B2 => gl_rom_rom_633(0), ZN => gl_rom_n_652);
  gl_rom_g35766 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_220(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_222(1), ZN => gl_rom_n_651);
  gl_rom_g35767 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_298(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_302(0), ZN => gl_rom_n_650);
  gl_rom_g35768 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_216(1), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_219(1), ZN => gl_rom_n_649);
  gl_rom_g35769 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_672(0), B1 => FE_OFN20_gl_rom_n_21, B2 => gl_rom_rom_673(0), ZN => gl_rom_n_648);
  gl_rom_g35770 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_226(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_231(1), ZN => gl_rom_n_647);
  gl_rom_g35771 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_228(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_230(1), ZN => gl_rom_n_646);
  gl_rom_g35772 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_21, A2 => gl_rom_rom_297(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_301(0), ZN => gl_rom_n_645);
  gl_rom_g35773 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_22, A2 => gl_rom_rom_229(1), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_227(1), ZN => gl_rom_n_644);
  gl_rom_g35774 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_296(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_299(0), ZN => gl_rom_n_643);
  gl_rom_g35775 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_224(1), B1 => FE_OFN23_gl_rom_n_21, B2 => gl_rom_rom_225(1), ZN => gl_rom_n_642);
  gl_rom_g35776 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_976(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_977(0), ZN => gl_rom_n_641);
  gl_rom_g35777 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_202(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_207(1), ZN => gl_rom_n_640);
  gl_rom_g35778 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_917(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_915(0), ZN => gl_rom_n_639);
  gl_rom_g35779 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_201(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_205(1), ZN => gl_rom_n_638);
  gl_rom_g35780 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_21, A2 => gl_rom_rom_281(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_285(0), ZN => gl_rom_n_637);
  gl_rom_g35781 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_912(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_913(0), ZN => gl_rom_n_636);
  gl_rom_g35782 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_204(1), B1 => FE_OFN4_gl_rom_n_16, B2 => gl_rom_rom_206(1), ZN => gl_rom_n_635);
  gl_rom_g35783 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_200(1), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_203(1), ZN => gl_rom_n_634);
  gl_rom_g35784 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_284(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_286(0), ZN => gl_rom_n_633);
  gl_rom_g35785 : AOI22D0BWP7T port map(A1 => FE_OFN3_gl_rom_n_16, A2 => gl_rom_rom_694(0), B1 => FE_OFN11_gl_rom_n_22, B2 => gl_rom_rom_693(0), ZN => gl_rom_n_632);
  gl_rom_g35786 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_193(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_197(1), ZN => gl_rom_n_631);
  gl_rom_g35787 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_282(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_283(0), ZN => gl_rom_n_630);
  gl_rom_g35788 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_196(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_198(1), ZN => gl_rom_n_629);
  gl_rom_g35789 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_617(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_621(0), ZN => gl_rom_n_628);
  gl_rom_g35790 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_280(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_287(0), ZN => gl_rom_n_627);
  gl_rom_g35791 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_194(1), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_195(1), ZN => gl_rom_n_626);
  gl_rom_g35792 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_192(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_199(1), ZN => gl_rom_n_625);
  gl_rom_g35793 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_692(0), B1 => FE_OFN19_gl_rom_n_21, B2 => gl_rom_rom_689(0), ZN => gl_rom_n_624);
  gl_rom_g35794 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_620(0), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_622(0), ZN => gl_rom_n_623);
  gl_rom_g35795 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_316(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_319(1), ZN => gl_rom_n_622);
  gl_rom_g35796 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_21, A2 => gl_rom_rom_289(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_293(0), ZN => gl_rom_n_621);
  gl_rom_g35797 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_314(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_318(1), ZN => gl_rom_n_620);
  gl_rom_g35798 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_690(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_695(0), ZN => gl_rom_n_619);
  gl_rom_g35799 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_292(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_294(0), ZN => gl_rom_n_618);
  gl_rom_g35800 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_313(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_317(1), ZN => gl_rom_n_617);
  gl_rom_g35801 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_688(0), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_691(0), ZN => gl_rom_n_616);
  gl_rom_g35802 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_312(1), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_315(1), ZN => gl_rom_n_615);
  gl_rom_g35803 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_290(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_291(0), ZN => gl_rom_n_614);
  gl_rom_g35804 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_300(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_303(1), ZN => gl_rom_n_613);
  gl_rom_g35805 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_298(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_302(1), ZN => gl_rom_n_612);
  gl_rom_g35806 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_297(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_301(1), ZN => gl_rom_n_611);
  gl_rom_g35807 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_296(1), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_299(1), ZN => gl_rom_n_610);
  gl_rom_g35808 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_288(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_295(0), ZN => gl_rom_n_609);
  gl_rom_g35809 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_618(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_619(0), ZN => gl_rom_n_608);
  gl_rom_g35810 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_308(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_311(1), ZN => gl_rom_n_607);
  gl_rom_g35811 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_306(1), B1 => FE_OFN4_gl_rom_n_16, B2 => gl_rom_rom_310(1), ZN => gl_rom_n_606);
  gl_rom_g35812 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_306(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_311(0), ZN => gl_rom_n_605);
  gl_rom_g35813 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_1001(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_1005(0), ZN => gl_rom_n_604);
  gl_rom_g35814 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_305(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_309(1), ZN => gl_rom_n_603);
  gl_rom_g35815 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_304(1), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_307(1), ZN => gl_rom_n_602);
  gl_rom_g35816 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_308(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_310(0), ZN => gl_rom_n_601);
  gl_rom_g35817 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_658(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_663(0), ZN => gl_rom_n_600);
  gl_rom_g35818 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_274(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_279(1), ZN => gl_rom_n_599);
  gl_rom_g35819 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_22, A2 => gl_rom_rom_309(0), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_307(0), ZN => gl_rom_n_598);
  gl_rom_g35820 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_273(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_277(1), ZN => gl_rom_n_597);
  gl_rom_g35821 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_21, A2 => gl_rom_rom_657(0), B1 => FE_OFN11_gl_rom_n_22, B2 => gl_rom_rom_661(0), ZN => gl_rom_n_596);
  gl_rom_g35822 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_276(1), B1 => FE_OFN4_gl_rom_n_16, B2 => gl_rom_rom_278(1), ZN => gl_rom_n_595);
  gl_rom_g35823 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_272(1), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_275(1), ZN => gl_rom_n_594);
  gl_rom_g35824 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_304(0), B1 => FE_OFN19_gl_rom_n_21, B2 => gl_rom_rom_305(0), ZN => gl_rom_n_593);
  gl_rom_g35825 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_282(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_287(1), ZN => gl_rom_n_592);
  gl_rom_g35826 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_274(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_279(0), ZN => gl_rom_n_591);
  gl_rom_g35827 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_281(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_285(1), ZN => gl_rom_n_590);
  gl_rom_g35828 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_616(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_623(0), ZN => gl_rom_n_589);
  gl_rom_g35829 : AOI22D0BWP7T port map(A1 => FE_OFN1_gl_rom_n_16, A2 => gl_rom_rom_662(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_659(0), ZN => gl_rom_n_588);
  gl_rom_g35830 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_284(1), B1 => FE_OFN4_gl_rom_n_16, B2 => gl_rom_rom_286(1), ZN => gl_rom_n_587);
  gl_rom_g35831 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_280(1), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_283(1), ZN => gl_rom_n_586);
  gl_rom_g35832 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_21, A2 => gl_rom_rom_273(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_277(0), ZN => gl_rom_n_585);
  gl_rom_g35833 : AOI22D0BWP7T port map(A1 => FE_OFN3_gl_rom_n_16, A2 => gl_rom_rom_278(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_275(0), ZN => gl_rom_n_584);
  gl_rom_g35834 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_290(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_295(1), ZN => gl_rom_n_583);
  gl_rom_g35835 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_289(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_293(1), ZN => gl_rom_n_582);
  gl_rom_g35836 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_656(0), B1 => FE_OFN7_gl_rom_n_18, B2 => gl_rom_rom_660(0), ZN => gl_rom_n_581);
  gl_rom_g35837 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_292(1), B1 => FE_OFN4_gl_rom_n_16, B2 => gl_rom_rom_294(1), ZN => gl_rom_n_580);
  gl_rom_g35838 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_272(0), B1 => FE_OFN7_gl_rom_n_18, B2 => gl_rom_rom_276(0), ZN => gl_rom_n_579);
  gl_rom_g35839 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_288(1), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_291(1), ZN => gl_rom_n_578);
  gl_rom_g35840 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_1004(0), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_1006(0), ZN => gl_rom_n_577);
  gl_rom_g35841 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_268(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_271(1), ZN => gl_rom_n_576);
  gl_rom_g35842 : AOI22D0BWP7T port map(A1 => FE_OFN0_gl_rom_n_16, A2 => gl_rom_rom_926(0), B1 => FE_OFN11_gl_rom_n_22, B2 => gl_rom_rom_925(0), ZN => gl_rom_n_575);
  gl_rom_g35843 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_266(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_271(0), ZN => gl_rom_n_574);
  gl_rom_g35844 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_266(1), B1 => FE_OFN4_gl_rom_n_16, B2 => gl_rom_rom_270(1), ZN => gl_rom_n_573);
  gl_rom_g35845 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_265(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_269(1), ZN => gl_rom_n_572);
  gl_rom_g35846 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_652(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_655(0), ZN => gl_rom_n_571);
  gl_rom_g35847 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_268(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_270(0), ZN => gl_rom_n_570);
  gl_rom_g35848 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_264(1), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_267(1), ZN => gl_rom_n_569);
  gl_rom_g35849 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_602(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_607(0), ZN => gl_rom_n_568);
  gl_rom_g35850 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_258(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_263(1), ZN => gl_rom_n_567);
  gl_rom_g35851 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_22, A2 => gl_rom_rom_269(0), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_267(0), ZN => gl_rom_n_566);
  gl_rom_g35852 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_257(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_261(1), ZN => gl_rom_n_565);
  gl_rom_g35853 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_264(0), B1 => FE_OFN19_gl_rom_n_21, B2 => gl_rom_rom_265(0), ZN => gl_rom_n_564);
  gl_rom_g35854 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_260(1), B1 => FE_OFN4_gl_rom_n_16, B2 => gl_rom_rom_262(1), ZN => gl_rom_n_563);
  gl_rom_g35855 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_256(1), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_259(1), ZN => gl_rom_n_562);
  gl_rom_g35856 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_650(0), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_654(0), ZN => gl_rom_n_561);
  gl_rom_g35857 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_258(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_263(0), ZN => gl_rom_n_560);
  gl_rom_g35858 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_346(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_351(1), ZN => gl_rom_n_559);
  gl_rom_g35859 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_604(0), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_606(0), ZN => gl_rom_n_558);
  gl_rom_g35860 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_21, A2 => gl_rom_rom_345(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_349(1), ZN => gl_rom_n_557);
  gl_rom_g35861 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_21, A2 => gl_rom_rom_257(0), B1 => FE_OFN11_gl_rom_n_22, B2 => gl_rom_rom_261(0), ZN => gl_rom_n_556);
  gl_rom_g35862 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_348(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_350(1), ZN => gl_rom_n_555);
  gl_rom_g35863 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_21, A2 => gl_rom_rom_649(0), B1 => FE_OFN11_gl_rom_n_22, B2 => gl_rom_rom_653(0), ZN => gl_rom_n_554);
  gl_rom_g35864 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_344(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_347(1), ZN => gl_rom_n_553);
  gl_rom_g35865 : AOI22D0BWP7T port map(A1 => FE_OFN3_gl_rom_n_16, A2 => gl_rom_rom_262(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_259(0), ZN => gl_rom_n_552);
  gl_rom_g35866 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_648(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_651(0), ZN => gl_rom_n_551);
  gl_rom_g35867 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_890(1), B1 => FE_OFN4_gl_rom_n_16, B2 => gl_rom_rom_894(1), ZN => gl_rom_n_550);
  gl_rom_g35868 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_356(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_358(1), ZN => gl_rom_n_549);
  gl_rom_g35869 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_256(0), B1 => FE_OFN7_gl_rom_n_18, B2 => gl_rom_rom_260(0), ZN => gl_rom_n_548);
  gl_rom_g35870 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_354(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_355(1), ZN => gl_rom_n_547);
  gl_rom_g35871 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_352(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_359(1), ZN => gl_rom_n_546);
  gl_rom_g35872 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_924(0), B1 => FE_OFN20_gl_rom_n_21, B2 => gl_rom_rom_921(0), ZN => gl_rom_n_545);
  gl_rom_g35873 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_370(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_375(1), ZN => gl_rom_n_544);
  gl_rom_g35874 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_369(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_373(1), ZN => gl_rom_n_543);
  gl_rom_g35875 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_22, A2 => gl_rom_rom_605(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_603(0), ZN => gl_rom_n_542);
  gl_rom_g35876 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_188(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_191(0), ZN => gl_rom_n_541);
  gl_rom_g35877 : AOI22D0BWP7T port map(A1 => FE_OFN3_gl_rom_n_16, A2 => gl_rom_rom_646(0), B1 => FE_OFN11_gl_rom_n_22, B2 => gl_rom_rom_645(0), ZN => gl_rom_n_540);
  gl_rom_g35878 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_372(1), B1 => FE_OFN4_gl_rom_n_16, B2 => gl_rom_rom_374(1), ZN => gl_rom_n_539);
  gl_rom_g35879 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_186(0), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_190(0), ZN => gl_rom_n_538);
  gl_rom_g35880 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_368(1), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_371(1), ZN => gl_rom_n_537);
  gl_rom_g35881 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_338(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_343(1), ZN => gl_rom_n_536);
  gl_rom_g35882 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_185(0), B1 => FE_OFN11_gl_rom_n_22, B2 => gl_rom_rom_189(0), ZN => gl_rom_n_535);
  gl_rom_g35883 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_337(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_341(1), ZN => gl_rom_n_534);
  gl_rom_g35884 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_644(0), B1 => FE_OFN19_gl_rom_n_21, B2 => gl_rom_rom_641(0), ZN => gl_rom_n_533);
  gl_rom_g35885 : AOI22D0BWP7T port map(A1 => FE_OFN4_gl_rom_n_16, A2 => gl_rom_rom_342(1), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_339(1), ZN => gl_rom_n_532);
  gl_rom_g35886 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_184(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_187(0), ZN => gl_rom_n_531);
  gl_rom_g35887 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_336(1), B1 => FE_OFN7_gl_rom_n_18, B2 => gl_rom_rom_340(1), ZN => gl_rom_n_530);
  gl_rom_g35888 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_600(0), B1 => FE_OFN20_gl_rom_n_21, B2 => gl_rom_rom_601(0), ZN => gl_rom_n_529);
  gl_rom_g35889 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_378(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_383(1), ZN => gl_rom_n_528);
  gl_rom_g35890 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_642(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_647(0), ZN => gl_rom_n_527);
  gl_rom_g35891 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_380(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_382(1), ZN => gl_rom_n_526);
  gl_rom_g35892 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_169(0), B1 => FE_OFN11_gl_rom_n_22, B2 => gl_rom_rom_173(0), ZN => gl_rom_n_525);
  gl_rom_g35893 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_172(0), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_174(0), ZN => gl_rom_n_524);
  gl_rom_g35894 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_22, A2 => gl_rom_rom_381(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_379(1), ZN => gl_rom_n_523);
  gl_rom_g35895 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_376(1), B1 => FE_OFN23_gl_rom_n_21, B2 => gl_rom_rom_377(1), ZN => gl_rom_n_522);
  gl_rom_g35896 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_362(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_367(1), ZN => gl_rom_n_521);
  gl_rom_g35897 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_640(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_643(0), ZN => gl_rom_n_520);
  gl_rom_g35898 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_170(0), B1 => FE_OFN17_gl_rom_n_15, B2 => gl_rom_rom_171(0), ZN => gl_rom_n_519);
  gl_rom_g35899 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_364(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_366(1), ZN => gl_rom_n_518);
  gl_rom_g35900 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_168(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_175(0), ZN => gl_rom_n_517);
  gl_rom_g35901 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_22, A2 => gl_rom_rom_365(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_363(1), ZN => gl_rom_n_516);
  gl_rom_g35902 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_360(1), B1 => FE_OFN23_gl_rom_n_21, B2 => gl_rom_rom_361(1), ZN => gl_rom_n_515);
  gl_rom_g35903 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_922(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_927(0), ZN => gl_rom_n_514);
  gl_rom_g35904 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_332(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_335(1), ZN => gl_rom_n_513);
  gl_rom_g35905 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_330(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_334(1), ZN => gl_rom_n_512);
  gl_rom_g35906 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_154(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_159(0), ZN => gl_rom_n_511);
  gl_rom_g35907 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_610(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_615(0), ZN => gl_rom_n_510);
  gl_rom_g35908 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_329(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_333(1), ZN => gl_rom_n_509);
  gl_rom_g35909 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_328(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_331(1), ZN => gl_rom_n_508);
  gl_rom_g35910 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_156(0), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_158(0), ZN => gl_rom_n_507);
  gl_rom_g35911 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_324(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_327(1), ZN => gl_rom_n_506);
  gl_rom_g35912 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_21, A2 => gl_rom_rom_561(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_565(0), ZN => gl_rom_n_505);
  gl_rom_g35913 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_22, A2 => gl_rom_rom_157(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_155(0), ZN => gl_rom_n_504);
  gl_rom_g35914 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_322(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_326(1), ZN => gl_rom_n_503);
  gl_rom_g35915 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_564(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_566(0), ZN => gl_rom_n_502);
  gl_rom_g35916 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_152(0), B1 => FE_OFN20_gl_rom_n_21, B2 => gl_rom_rom_153(0), ZN => gl_rom_n_501);
  gl_rom_g35917 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_321(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_325(1), ZN => gl_rom_n_500);
  gl_rom_g35918 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_320(1), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_323(1), ZN => gl_rom_n_499);
  gl_rom_g35919 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_609(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_613(0), ZN => gl_rom_n_498);
  gl_rom_g35920 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_122(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_127(1), ZN => gl_rom_n_497);
  gl_rom_g35921 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_164(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_167(0), ZN => gl_rom_n_496);
  gl_rom_g35922 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_121(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_125(1), ZN => gl_rom_n_495);
  gl_rom_g35923 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_124(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_126(1), ZN => gl_rom_n_494);
  gl_rom_g35924 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_562(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_563(0), ZN => gl_rom_n_493);
  gl_rom_g35925 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_162(0), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_166(0), ZN => gl_rom_n_492);
  gl_rom_g35926 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_120(1), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_123(1), ZN => gl_rom_n_491);
  gl_rom_g35927 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_920(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_923(0), ZN => gl_rom_n_490);
  gl_rom_g35928 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_108(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_111(1), ZN => gl_rom_n_489);
  gl_rom_g35929 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_161(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_165(0), ZN => gl_rom_n_488);
  gl_rom_g35930 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_560(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_567(0), ZN => gl_rom_n_487);
  gl_rom_g35931 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_106(1), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_110(1), ZN => gl_rom_n_486);
  gl_rom_g35932 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_160(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_163(0), ZN => gl_rom_n_485);
  gl_rom_g35933 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_105(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_109(1), ZN => gl_rom_n_484);
  gl_rom_g35934 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_104(1), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_107(1), ZN => gl_rom_n_483);
  gl_rom_g35935 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_1002(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_1003(0), ZN => gl_rom_n_482);
  gl_rom_g35936 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_92(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_95(1), ZN => gl_rom_n_481);
  gl_rom_g35937 : AOI22D0BWP7T port map(A1 => FE_OFN1_gl_rom_n_16, A2 => gl_rom_rom_614(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_611(0), ZN => gl_rom_n_480);
  gl_rom_g35938 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_90(1), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_94(1), ZN => gl_rom_n_479);
  gl_rom_g35939 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_178(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_183(0), ZN => gl_rom_n_478);
  gl_rom_g35940 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_89(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_93(1), ZN => gl_rom_n_477);
  gl_rom_g35941 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_608(0), B1 => FE_OFN6_gl_rom_n_18, B2 => gl_rom_rom_612(0), ZN => gl_rom_n_476);
  gl_rom_g35942 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_180(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_182(0), ZN => gl_rom_n_475);
  gl_rom_g35943 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_88(1), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_91(1), ZN => gl_rom_n_474);
  gl_rom_g35944 : AOI22D0BWP7T port map(A1 => FE_OFN3_gl_rom_n_16, A2 => gl_rom_rom_534(0), B1 => FE_OFN11_gl_rom_n_22, B2 => gl_rom_rom_533(0), ZN => gl_rom_n_473);
  gl_rom_g35945 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_97(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_101(1), ZN => gl_rom_n_472);
  gl_rom_g35946 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_532(0), B1 => FE_OFN19_gl_rom_n_21, B2 => gl_rom_rom_529(0), ZN => gl_rom_n_471);
  gl_rom_g35947 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_100(1), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_102(1), ZN => gl_rom_n_470);
  gl_rom_g35948 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_22, A2 => gl_rom_rom_181(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_179(0), ZN => gl_rom_n_469);
  gl_rom_g35949 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_98(1), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_99(1), ZN => gl_rom_n_468);
  gl_rom_g35950 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_176(0), B1 => FE_OFN19_gl_rom_n_21, B2 => gl_rom_rom_177(0), ZN => gl_rom_n_467);
  gl_rom_g35951 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_96(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_103(1), ZN => gl_rom_n_466);
  gl_rom_g35952 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_114(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_119(1), ZN => gl_rom_n_465);
  gl_rom_g35953 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_146(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_151(0), ZN => gl_rom_n_464);
  gl_rom_g35954 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_21, A2 => gl_rom_rom_113(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_117(1), ZN => gl_rom_n_463);
  gl_rom_g35955 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_530(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_535(0), ZN => gl_rom_n_462);
  gl_rom_g35956 : AOI22D0BWP7T port map(A1 => FE_OFN0_gl_rom_n_16, A2 => gl_rom_rom_118(1), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_115(1), ZN => gl_rom_n_461);
  gl_rom_g35957 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_148(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_150(0), ZN => gl_rom_n_460);
  gl_rom_g35958 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_112(1), B1 => FE_OFN5_gl_rom_n_18, B2 => gl_rom_rom_116(1), ZN => gl_rom_n_459);
  gl_rom_g35959 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_82(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_87(1), ZN => gl_rom_n_458);
  gl_rom_g35960 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_22, A2 => gl_rom_rom_149(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_147(0), ZN => gl_rom_n_457);
  gl_rom_g35961 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_84(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_86(1), ZN => gl_rom_n_456);
  gl_rom_g35962 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_1000(0), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_1007(0), ZN => gl_rom_n_455);
  gl_rom_g35963 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_528(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_531(0), ZN => gl_rom_n_454);
  gl_rom_g35964 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_85(1), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_83(1), ZN => gl_rom_n_453);
  gl_rom_g35965 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_144(0), B1 => FE_OFN19_gl_rom_n_21, B2 => gl_rom_rom_145(0), ZN => gl_rom_n_452);
  gl_rom_g35966 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_80(1), B1 => FE_OFN23_gl_rom_n_21, B2 => gl_rom_rom_81(1), ZN => gl_rom_n_451);
  gl_rom_g35967 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_930(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_935(0), ZN => gl_rom_n_450);
  gl_rom_g35968 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_73(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_77(1), ZN => gl_rom_n_449);
  gl_rom_g35969 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_138(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_143(0), ZN => gl_rom_n_448);
  gl_rom_g35970 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_76(1), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_78(1), ZN => gl_rom_n_447);
  gl_rom_g35971 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_74(1), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_75(1), ZN => gl_rom_n_446);
  gl_rom_g35972 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_625(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_629(0), ZN => gl_rom_n_445);
  gl_rom_g35973 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_140(0), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_142(0), ZN => gl_rom_n_444);
  gl_rom_g35974 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_72(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_79(1), ZN => gl_rom_n_443);
  gl_rom_g35975 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_538(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_543(0), ZN => gl_rom_n_442);
  gl_rom_g35976 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_68(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_71(1), ZN => gl_rom_n_441);
  gl_rom_g35977 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_22, A2 => gl_rom_rom_141(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_139(0), ZN => gl_rom_n_440);
  gl_rom_g35978 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_66(1), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_70(1), ZN => gl_rom_n_439);
  gl_rom_g35979 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_136(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_137(0), ZN => gl_rom_n_438);
  gl_rom_g35980 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_65(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_69(1), ZN => gl_rom_n_437);
  gl_rom_g35981 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_64(1), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_67(1), ZN => gl_rom_n_436);
  gl_rom_g35982 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_537(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_541(0), ZN => gl_rom_n_435);
  gl_rom_g35983 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_130(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_135(0), ZN => gl_rom_n_434);
  gl_rom_g35984 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_180(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_183(1), ZN => gl_rom_n_433);
  gl_rom_g35985 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_628(0), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_630(0), ZN => gl_rom_n_432);
  gl_rom_g35986 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_178(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_182(1), ZN => gl_rom_n_431);
  gl_rom_g35987 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_21, A2 => gl_rom_rom_129(0), B1 => FE_OFN11_gl_rom_n_22, B2 => gl_rom_rom_133(0), ZN => gl_rom_n_430);
  gl_rom_g35988 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_21, A2 => gl_rom_rom_177(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_181(1), ZN => gl_rom_n_429);
  gl_rom_g35989 : AOI22D0BWP7T port map(A1 => FE_OFN1_gl_rom_n_16, A2 => gl_rom_rom_542(0), B1 => FE_OFN17_gl_rom_n_15, B2 => gl_rom_rom_539(0), ZN => gl_rom_n_428);
  gl_rom_g35990 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_176(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_179(1), ZN => gl_rom_n_427);
  gl_rom_g35991 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_132(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_134(0), ZN => gl_rom_n_426);
  gl_rom_g35992 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_986(0), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_991(0), ZN => gl_rom_n_425);
  gl_rom_g35993 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_536(0), B1 => FE_OFN5_gl_rom_n_18, B2 => gl_rom_rom_540(0), ZN => gl_rom_n_424);
  gl_rom_g35994 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_148(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_151(1), ZN => gl_rom_n_423);
  gl_rom_g35995 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_146(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_150(1), ZN => gl_rom_n_422);
  gl_rom_g35996 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_128(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_131(0), ZN => gl_rom_n_421);
  gl_rom_g35997 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_21, A2 => gl_rom_rom_145(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_149(1), ZN => gl_rom_n_420);
  gl_rom_g35998 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_929(0), B1 => FE_OFN11_gl_rom_n_22, B2 => gl_rom_rom_933(0), ZN => gl_rom_n_419);
  gl_rom_g35999 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_144(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_147(1), ZN => gl_rom_n_418);
  gl_rom_g36000 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_156(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_159(1), ZN => gl_rom_n_417);
  gl_rom_g36001 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_626(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_627(0), ZN => gl_rom_n_416);
  gl_rom_g36002 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_154(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_158(1), ZN => gl_rom_n_415);
  gl_rom_g36003 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_58(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_63(0), ZN => gl_rom_n_414);
  gl_rom_g36004 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_153(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_157(1), ZN => gl_rom_n_413);
  gl_rom_g36005 : AOI22D0BWP7T port map(A1 => FE_OFN1_gl_rom_n_16, A2 => gl_rom_rom_550(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_549(0), ZN => gl_rom_n_412);
  gl_rom_g36006 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_152(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_155(1), ZN => gl_rom_n_411);
  gl_rom_g36007 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_57(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_61(0), ZN => gl_rom_n_410);
  gl_rom_g36008 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_162(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_167(1), ZN => gl_rom_n_409);
  gl_rom_g36009 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_164(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_166(1), ZN => gl_rom_n_408);
  gl_rom_g36010 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_60(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_62(0), ZN => gl_rom_n_407);
  gl_rom_g36011 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_56(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_59(0), ZN => gl_rom_n_406);
  gl_rom_g36012 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_22, A2 => gl_rom_rom_165(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_163(1), ZN => gl_rom_n_405);
  gl_rom_g36013 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_160(1), B1 => FE_OFN22_gl_rom_n_21, B2 => gl_rom_rom_161(1), ZN => gl_rom_n_404);
  gl_rom_g36014 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_548(0), B1 => FE_OFN20_gl_rom_n_21, B2 => gl_rom_rom_545(0), ZN => gl_rom_n_403);
  gl_rom_g36015 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_188(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_191(1), ZN => gl_rom_n_402);
  gl_rom_g36016 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_624(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_631(0), ZN => gl_rom_n_401);
  gl_rom_g36017 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_44(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_47(0), ZN => gl_rom_n_400);
  gl_rom_g36018 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_186(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_190(1), ZN => gl_rom_n_399);
  gl_rom_g36019 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_546(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_551(0), ZN => gl_rom_n_398);
  gl_rom_g36020 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_21, A2 => gl_rom_rom_185(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_189(1), ZN => gl_rom_n_397);
  gl_rom_g36021 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_42(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_46(0), ZN => gl_rom_n_396);
  gl_rom_g36022 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_184(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_187(1), ZN => gl_rom_n_395);
  gl_rom_g36023 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_170(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_175(1), ZN => gl_rom_n_394);
  gl_rom_g36024 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_544(0), B1 => FE_OFN17_gl_rom_n_15, B2 => gl_rom_rom_547(0), ZN => gl_rom_n_393);
  gl_rom_g36025 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_41(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_45(0), ZN => gl_rom_n_392);
  gl_rom_g36026 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_172(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_174(1), ZN => gl_rom_n_391);
  gl_rom_g36027 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_40(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_43(0), ZN => gl_rom_n_390);
  gl_rom_g36028 : AOI22D0BWP7T port map(A1 => FE_OFN12_gl_rom_n_22, A2 => gl_rom_rom_173(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_171(1), ZN => gl_rom_n_389);
  gl_rom_g36029 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_168(1), B1 => FE_OFN23_gl_rom_n_21, B2 => gl_rom_rom_169(1), ZN => gl_rom_n_388);
  gl_rom_g36030 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_1013(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_1011(0), ZN => gl_rom_n_387);
  gl_rom_g36031 : AOI22D0BWP7T port map(A1 => FE_OFN0_gl_rom_n_16, A2 => gl_rom_rom_934(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_931(0), ZN => gl_rom_n_386);
  gl_rom_g36032 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_140(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_143(1), ZN => gl_rom_n_385);
  gl_rom_g36033 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_594(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_599(0), ZN => gl_rom_n_384);
  gl_rom_g36034 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_138(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_142(1), ZN => gl_rom_n_383);
  gl_rom_g36035 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_50(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_55(0), ZN => gl_rom_n_382);
  gl_rom_g36036 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_137(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_141(1), ZN => gl_rom_n_381);
  gl_rom_g36037 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_52(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_54(0), ZN => gl_rom_n_380);
  gl_rom_g36038 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_136(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_139(1), ZN => gl_rom_n_379);
  gl_rom_g36039 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_570(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_575(0), ZN => gl_rom_n_378);
  gl_rom_g36040 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_132(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_135(1), ZN => gl_rom_n_377);
  gl_rom_g36041 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_22, A2 => gl_rom_rom_53(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_51(0), ZN => gl_rom_n_376);
  gl_rom_g36042 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_130(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_134(1), ZN => gl_rom_n_375);
  gl_rom_g36043 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_572(0), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_574(0), ZN => gl_rom_n_374);
  gl_rom_g36044 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_48(0), B1 => FE_OFN20_gl_rom_n_21, B2 => gl_rom_rom_49(0), ZN => gl_rom_n_373);
  gl_rom_g36045 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_129(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_133(1), ZN => gl_rom_n_372);
  gl_rom_g36046 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_128(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_131(1), ZN => gl_rom_n_371);
  gl_rom_g36047 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_593(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_597(0), ZN => gl_rom_n_370);
  gl_rom_g36048 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_60(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_63(1), ZN => gl_rom_n_369);
  gl_rom_g36049 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_17(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_21(0), ZN => gl_rom_n_368);
  gl_rom_g36050 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_58(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_62(1), ZN => gl_rom_n_367);
  gl_rom_g36051 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_57(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_61(1), ZN => gl_rom_n_366);
  gl_rom_g36052 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_20(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_22(0), ZN => gl_rom_n_365);
  gl_rom_g36053 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_56(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_59(1), ZN => gl_rom_n_364);
  gl_rom_g36054 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_928(0), B1 => FE_OFN5_gl_rom_n_18, B2 => gl_rom_rom_932(0), ZN => gl_rom_n_363);
  gl_rom_g36055 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_22, A2 => gl_rom_rom_573(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_571(0), ZN => gl_rom_n_362);
  gl_rom_g36056 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_18(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_19(0), ZN => gl_rom_n_361);
  gl_rom_g36057 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_44(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_47(1), ZN => gl_rom_n_360);
  gl_rom_g36058 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_568(0), B1 => FE_OFN20_gl_rom_n_21, B2 => gl_rom_rom_569(0), ZN => gl_rom_n_359);
  gl_rom_g36059 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_42(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_46(1), ZN => gl_rom_n_358);
  gl_rom_g36060 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_16(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_23(0), ZN => gl_rom_n_357);
  gl_rom_g36061 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_41(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_45(1), ZN => gl_rom_n_356);
  gl_rom_g36062 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_40(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_43(1), ZN => gl_rom_n_355);
  gl_rom_g36063 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_52(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_55(1), ZN => gl_rom_n_354);
  gl_rom_g36064 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_596(0), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_598(0), ZN => gl_rom_n_353);
  gl_rom_g36065 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_26(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_31(0), ZN => gl_rom_n_352);
  gl_rom_g36066 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_50(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_54(1), ZN => gl_rom_n_351);
  gl_rom_g36067 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_553(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_557(0), ZN => gl_rom_n_350);
  gl_rom_g36068 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_49(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_53(1), ZN => gl_rom_n_349);
  gl_rom_g36069 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_25(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_29(0), ZN => gl_rom_n_348);
  gl_rom_g36070 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_48(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_51(1), ZN => gl_rom_n_347);
  gl_rom_g36071 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_17(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_21(1), ZN => gl_rom_n_346);
  gl_rom_g36072 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_969(0), B1 => FE_OFN11_gl_rom_n_22, B2 => gl_rom_rom_973(0), ZN => gl_rom_n_345);
  gl_rom_g36073 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_20(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_22(1), ZN => gl_rom_n_344);
  gl_rom_g36074 : AOI22D0BWP7T port map(A1 => FE_OFN3_gl_rom_n_16, A2 => gl_rom_rom_30(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_27(0), ZN => gl_rom_n_343);
  gl_rom_g36075 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_592(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_595(0), ZN => gl_rom_n_342);
  gl_rom_g36076 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_556(0), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_558(0), ZN => gl_rom_n_341);
  gl_rom_g36077 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_18(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_19(1), ZN => gl_rom_n_340);
  gl_rom_g36078 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_24(0), B1 => FE_OFN6_gl_rom_n_18, B2 => gl_rom_rom_28(0), ZN => gl_rom_n_339);
  gl_rom_g36079 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_16(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_23(1), ZN => gl_rom_n_338);
  gl_rom_g36080 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_28(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_31(1), ZN => gl_rom_n_337);
  gl_rom_g36081 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_34(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_39(0), ZN => gl_rom_n_336);
  gl_rom_g36082 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_26(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_30(1), ZN => gl_rom_n_335);
  gl_rom_g36083 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_36(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_38(0), ZN => gl_rom_n_334);
  gl_rom_g36084 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_25(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_29(1), ZN => gl_rom_n_333);
  gl_rom_g36085 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_24(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_27(1), ZN => gl_rom_n_332);
  gl_rom_g36086 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_554(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_555(0), ZN => gl_rom_n_331);
  gl_rom_g36087 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_34(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_39(1), ZN => gl_rom_n_330);
  gl_rom_g36088 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_552(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_559(0), ZN => gl_rom_n_329);
  gl_rom_g36089 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_22, A2 => gl_rom_rom_37(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_35(0), ZN => gl_rom_n_328);
  gl_rom_g36090 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_33(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_37(1), ZN => gl_rom_n_327);
  gl_rom_g36091 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_988(0), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_990(0), ZN => gl_rom_n_326);
  gl_rom_g36092 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_32(0), B1 => FE_OFN20_gl_rom_n_21, B2 => gl_rom_rom_33(0), ZN => gl_rom_n_325);
  gl_rom_g36093 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_36(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_38(1), ZN => gl_rom_n_324);
  gl_rom_g36094 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_32(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_35(1), ZN => gl_rom_n_323);
  gl_rom_g36095 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_908(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_911(0), ZN => gl_rom_n_322);
  gl_rom_g36096 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_9(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_13(1), ZN => gl_rom_n_321);
  gl_rom_g36097 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_12(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_15(0), ZN => gl_rom_n_320);
  gl_rom_g36098 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_12(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_14(1), ZN => gl_rom_n_319);
  gl_rom_g36099 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_10(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_11(1), ZN => gl_rom_n_318);
  gl_rom_g36100 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_586(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_591(0), ZN => gl_rom_n_317);
  gl_rom_g36101 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_10(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_14(0), ZN => gl_rom_n_316);
  gl_rom_g36102 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_8(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_15(1), ZN => gl_rom_n_315);
  gl_rom_g36103 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_524(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_527(0), ZN => gl_rom_n_314);
  gl_rom_g36104 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_522(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_526(0), ZN => gl_rom_n_313);
  gl_rom_g36105 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_21, A2 => gl_rom_rom_9(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_13(0), ZN => gl_rom_n_312);
  gl_rom_g36106 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_2(1), B1 => gl_rom_n_17, B2 => gl_rom_rom_7(1), ZN => gl_rom_n_311);
  gl_rom_g36107 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_1(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_5(1), ZN => gl_rom_n_310);
  gl_rom_g36108 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_588(0), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_590(0), ZN => gl_rom_n_309);
  gl_rom_g36109 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_8(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_11(0), ZN => gl_rom_n_308);
  gl_rom_g36110 : AOI22D0BWP7T port map(A1 => gl_rom_n_18, A2 => gl_rom_rom_4(1), B1 => gl_rom_n_16, B2 => gl_rom_rom_6(1), ZN => gl_rom_n_307);
  gl_rom_g36111 : AOI22D0BWP7T port map(A1 => gl_rom_n_19, A2 => gl_rom_rom_0(1), B1 => gl_rom_n_15, B2 => gl_rom_rom_3(1), ZN => gl_rom_n_306);
  gl_rom_g36112 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_1(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_5(0), ZN => gl_rom_n_305);
  gl_rom_g36113 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_21, A2 => gl_rom_rom_521(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_525(0), ZN => gl_rom_n_304);
  gl_rom_g36114 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_4(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_6(0), ZN => gl_rom_n_303);
  gl_rom_g36115 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_906(0), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_910(0), ZN => gl_rom_n_302);
  gl_rom_g36116 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_520(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_523(0), ZN => gl_rom_n_301);
  gl_rom_g36117 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_2(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_3(0), ZN => gl_rom_n_300);
  gl_rom_g36118 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_0(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_7(0), ZN => gl_rom_n_299);
  gl_rom_g36119 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_22, A2 => gl_rom_rom_589(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_587(0), ZN => gl_rom_n_298);
  gl_rom_g36120 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_21, A2 => gl_rom_rom_513(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_517(0), ZN => gl_rom_n_297);
  gl_rom_g36121 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_516(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_518(0), ZN => gl_rom_n_296);
  gl_rom_g36122 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_892(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_895(1), ZN => gl_rom_n_295);
  gl_rom_g36123 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_21, A2 => gl_rom_rom_353(1), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_357(1), ZN => gl_rom_n_294);
  gl_rom_g36124 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_584(0), B1 => FE_OFN20_gl_rom_n_21, B2 => gl_rom_rom_585(0), ZN => gl_rom_n_293);
  gl_rom_g36125 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_889(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_893(1), ZN => gl_rom_n_292);
  gl_rom_g36126 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_514(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_515(0), ZN => gl_rom_n_291);
  gl_rom_g36127 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_888(1), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_891(1), ZN => gl_rom_n_290);
  gl_rom_g36128 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_972(0), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_974(0), ZN => gl_rom_n_289);
  gl_rom_g36129 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_905(0), B1 => FE_OFN11_gl_rom_n_22, B2 => gl_rom_rom_909(0), ZN => gl_rom_n_288);
  gl_rom_g36130 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_876(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_879(1), ZN => gl_rom_n_287);
  gl_rom_g36131 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_512(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_519(0), ZN => gl_rom_n_286);
  gl_rom_g36132 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_874(1), B1 => FE_OFN4_gl_rom_n_16, B2 => gl_rom_rom_878(1), ZN => gl_rom_n_285);
  gl_rom_g36133 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_873(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_877(1), ZN => gl_rom_n_284);
  gl_rom_g36134 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_872(1), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_875(1), ZN => gl_rom_n_283);
  gl_rom_g36135 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_578(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_583(0), ZN => gl_rom_n_282);
  gl_rom_g36136 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_580(0), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_582(0), ZN => gl_rom_n_281);
  gl_rom_g36137 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_860(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_863(1), ZN => gl_rom_n_280);
  gl_rom_g36138 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_904(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_907(0), ZN => gl_rom_n_279);
  gl_rom_g36139 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_858(1), B1 => FE_OFN4_gl_rom_n_16, B2 => gl_rom_rom_862(1), ZN => gl_rom_n_278);
  gl_rom_g36140 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_506(0), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_511(0), ZN => gl_rom_n_277);
  gl_rom_g36141 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_857(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_861(1), ZN => gl_rom_n_276);
  gl_rom_g36142 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_21, A2 => gl_rom_rom_505(0), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_509(0), ZN => gl_rom_n_275);
  gl_rom_g36143 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_856(1), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_859(1), ZN => gl_rom_n_274);
  gl_rom_g36144 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_868(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_871(1), ZN => gl_rom_n_273);
  gl_rom_g36145 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_866(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_870(1), ZN => gl_rom_n_272);
  gl_rom_g36146 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_989(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_987(0), ZN => gl_rom_n_271);
  gl_rom_g36147 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_22, A2 => gl_rom_rom_581(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_579(0), ZN => gl_rom_n_270);
  gl_rom_g36148 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_508(0), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_510(0), ZN => gl_rom_n_269);
  gl_rom_g36149 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_865(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_869(1), ZN => gl_rom_n_268);
  gl_rom_g36150 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_864(1), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_867(1), ZN => gl_rom_n_267);
  gl_rom_g36151 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_504(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_507(0), ZN => gl_rom_n_266);
  gl_rom_g36152 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_970(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_971(0), ZN => gl_rom_n_265);
  gl_rom_g36153 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_884(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_887(1), ZN => gl_rom_n_264);
  gl_rom_g36154 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_882(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_886(1), ZN => gl_rom_n_263);
  gl_rom_g36155 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_576(0), B1 => FE_OFN20_gl_rom_n_21, B2 => gl_rom_rom_577(0), ZN => gl_rom_n_262);
  gl_rom_g36156 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_492(0), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_495(0), ZN => gl_rom_n_261);
  gl_rom_g36157 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_881(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_885(1), ZN => gl_rom_n_260);
  gl_rom_g36158 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_490(0), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_494(0), ZN => gl_rom_n_259);
  gl_rom_g36159 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_880(1), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_883(1), ZN => gl_rom_n_258);
  gl_rom_g36160 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_968(0), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_975(0), ZN => gl_rom_n_257);
  gl_rom_g36161 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_852(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_855(1), ZN => gl_rom_n_256);
  gl_rom_g36162 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_850(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_854(1), ZN => gl_rom_n_255);
  gl_rom_g36163 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_21, A2 => gl_rom_rom_489(0), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_493(0), ZN => gl_rom_n_254);
  gl_rom_g36164 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_897(0), B1 => FE_OFN11_gl_rom_n_22, B2 => gl_rom_rom_901(0), ZN => gl_rom_n_253);
  gl_rom_g36165 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_849(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_853(1), ZN => gl_rom_n_252);
  gl_rom_g36166 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_848(1), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_851(1), ZN => gl_rom_n_251);
  gl_rom_g36167 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_488(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_491(0), ZN => gl_rom_n_250);
  gl_rom_g36168 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_900(0), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_902(0), ZN => gl_rom_n_249);
  gl_rom_g36169 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_841(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_845(1), ZN => gl_rom_n_248);
  gl_rom_g36170 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_844(1), B1 => FE_OFN4_gl_rom_n_16, B2 => gl_rom_rom_846(1), ZN => gl_rom_n_247);
  gl_rom_g36171 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_476(0), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_479(0), ZN => gl_rom_n_246);
  gl_rom_g36172 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_842(1), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_843(1), ZN => gl_rom_n_245);
  gl_rom_g36173 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_754(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_759(0), ZN => gl_rom_n_244);
  gl_rom_g36174 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_840(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_847(1), ZN => gl_rom_n_243);
  gl_rom_g36175 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_474(0), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_478(0), ZN => gl_rom_n_242);
  gl_rom_g36176 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_833(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_837(1), ZN => gl_rom_n_241);
  gl_rom_g36177 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_836(1), B1 => FE_OFN4_gl_rom_n_16, B2 => gl_rom_rom_838(1), ZN => gl_rom_n_240);
  gl_rom_g36178 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_473(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_477(0), ZN => gl_rom_n_239);
  gl_rom_g36179 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_834(1), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_835(1), ZN => gl_rom_n_238);
  gl_rom_g36180 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_472(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_475(0), ZN => gl_rom_n_237);
  gl_rom_g36181 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_832(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_839(1), ZN => gl_rom_n_236);
  gl_rom_g36182 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_21, A2 => gl_rom_rom_753(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_757(0), ZN => gl_rom_n_235);
  gl_rom_g36183 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_601(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_605(1), ZN => gl_rom_n_234);
  gl_rom_g36184 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_604(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_606(1), ZN => gl_rom_n_233);
  gl_rom_g36185 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_482(0), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_487(0), ZN => gl_rom_n_232);
  gl_rom_g36186 : AOI22D0BWP7T port map(A1 => FE_OFN3_gl_rom_n_16, A2 => gl_rom_rom_758(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_755(0), ZN => gl_rom_n_231);
  gl_rom_g36187 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_602(1), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_603(1), ZN => gl_rom_n_230);
  gl_rom_g36188 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_600(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_607(1), ZN => gl_rom_n_229);
  gl_rom_g36189 : AOI22D0BWP7T port map(A1 => FE_OFN23_gl_rom_n_21, A2 => gl_rom_rom_481(0), B1 => FE_OFN12_gl_rom_n_22, B2 => gl_rom_rom_485(0), ZN => gl_rom_n_228);
  gl_rom_g36190 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_752(0), B1 => FE_OFN6_gl_rom_n_18, B2 => gl_rom_rom_756(0), ZN => gl_rom_n_227);
  gl_rom_g36191 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_609(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_613(1), ZN => gl_rom_n_226);
  gl_rom_g36192 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_484(0), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_486(0), ZN => gl_rom_n_225);
  gl_rom_g36193 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_612(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_614(1), ZN => gl_rom_n_224);
  gl_rom_g36194 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_898(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_899(0), ZN => gl_rom_n_223);
  gl_rom_g36195 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_480(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_483(0), ZN => gl_rom_n_222);
  gl_rom_g36196 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_610(1), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_611(1), ZN => gl_rom_n_221);
  gl_rom_g36197 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_608(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_615(1), ZN => gl_rom_n_220);
  gl_rom_g36198 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_626(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_631(1), ZN => gl_rom_n_219);
  gl_rom_g36199 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_896(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_903(0), ZN => gl_rom_n_218);
  gl_rom_g36200 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_625(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_629(1), ZN => gl_rom_n_217);
  gl_rom_g36201 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_722(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_727(0), ZN => gl_rom_n_216);
  gl_rom_g36202 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_500(0), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_503(0), ZN => gl_rom_n_215);
  gl_rom_g36203 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_628(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_630(1), ZN => gl_rom_n_214);
  gl_rom_g36204 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_624(1), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_627(1), ZN => gl_rom_n_213);
  gl_rom_g36205 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_498(0), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_502(0), ZN => gl_rom_n_212);
  gl_rom_g36206 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_724(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_726(0), ZN => gl_rom_n_211);
  gl_rom_g36207 : AOI22D0BWP7T port map(A1 => FE_OFN0_gl_rom_n_16, A2 => gl_rom_rom_598(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_597(1), ZN => gl_rom_n_210);
  gl_rom_g36208 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_596(1), B1 => gl_rom_n_21, B2 => gl_rom_rom_593(1), ZN => gl_rom_n_209);
  gl_rom_g36209 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_497(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_501(0), ZN => gl_rom_n_208);
  gl_rom_g36210 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_594(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_599(1), ZN => gl_rom_n_207);
  gl_rom_g36211 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_592(1), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_595(1), ZN => gl_rom_n_206);
  gl_rom_g36212 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_496(0), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_499(0), ZN => gl_rom_n_205);
  gl_rom_g36213 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_634(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_639(1), ZN => gl_rom_n_204);
  gl_rom_g36214 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_984(0), B1 => FE_OFN20_gl_rom_n_21, B2 => gl_rom_rom_985(0), ZN => gl_rom_n_203);
  gl_rom_g36215 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_1008(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_1009(0), ZN => gl_rom_n_202);
  gl_rom_g36216 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_465(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_469(0), ZN => gl_rom_n_201);
  gl_rom_g36217 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_636(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_638(1), ZN => gl_rom_n_200);
  gl_rom_g36218 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_22, A2 => gl_rom_rom_725(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_723(0), ZN => gl_rom_n_199);
  gl_rom_g36219 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_637(1), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_635(1), ZN => gl_rom_n_198);
  gl_rom_g36220 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_468(0), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_470(0), ZN => gl_rom_n_197);
  gl_rom_g36221 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_632(1), B1 => gl_rom_n_21, B2 => gl_rom_rom_633(1), ZN => gl_rom_n_196);
  gl_rom_g36222 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_962(0), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_967(0), ZN => gl_rom_n_195);
  gl_rom_g36223 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_618(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_623(1), ZN => gl_rom_n_194);
  gl_rom_g36224 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_720(0), B1 => FE_OFN19_gl_rom_n_21, B2 => gl_rom_rom_721(0), ZN => gl_rom_n_193);
  gl_rom_g36225 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_617(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_621(1), ZN => gl_rom_n_192);
  gl_rom_g36226 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_466(0), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_467(0), ZN => gl_rom_n_191);
  gl_rom_g36227 : AOI22D0BWP7T port map(A1 => FE_OFN0_gl_rom_n_16, A2 => gl_rom_rom_622(1), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_619(1), ZN => gl_rom_n_190);
  gl_rom_g36228 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_464(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_471(0), ZN => gl_rom_n_189);
  gl_rom_g36229 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_616(1), B1 => FE_OFN5_gl_rom_n_18, B2 => gl_rom_rom_620(1), ZN => gl_rom_n_188);
  gl_rom_g36230 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_588(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_591(1), ZN => gl_rom_n_187);
  gl_rom_g36231 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_586(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_590(1), ZN => gl_rom_n_186);
  gl_rom_g36232 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_460(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_463(0), ZN => gl_rom_n_185);
  gl_rom_g36233 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_585(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_589(1), ZN => gl_rom_n_184);
  gl_rom_g36234 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_730(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_735(0), ZN => gl_rom_n_183);
  gl_rom_g36235 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_458(0), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_462(0), ZN => gl_rom_n_182);
  gl_rom_g36236 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_584(1), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_587(1), ZN => gl_rom_n_181);
  gl_rom_g36237 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_964(0), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_966(0), ZN => gl_rom_n_180);
  gl_rom_g36238 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_577(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_581(1), ZN => gl_rom_n_179);
  gl_rom_g36239 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_21, A2 => gl_rom_rom_729(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_733(0), ZN => gl_rom_n_178);
  gl_rom_g36240 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_580(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_582(1), ZN => gl_rom_n_177);
  gl_rom_g36241 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_457(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_461(0), ZN => gl_rom_n_176);
  gl_rom_g36242 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_857(0), B1 => FE_OFN11_gl_rom_n_22, B2 => gl_rom_rom_861(0), ZN => gl_rom_n_175);
  gl_rom_g36243 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_578(1), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_579(1), ZN => gl_rom_n_174);
  gl_rom_g36244 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_576(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_583(1), ZN => gl_rom_n_173);
  gl_rom_g36245 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_456(0), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_459(0), ZN => gl_rom_n_172);
  gl_rom_g36246 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_860(0), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_862(0), ZN => gl_rom_n_171);
  gl_rom_g36247 : AOI22D0BWP7T port map(A1 => FE_OFN4_gl_rom_n_16, A2 => gl_rom_rom_766(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_765(1), ZN => gl_rom_n_170);
  gl_rom_g36248 : AOI22D0BWP7T port map(A1 => FE_OFN3_gl_rom_n_16, A2 => gl_rom_rom_734(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_731(0), ZN => gl_rom_n_169);
  gl_rom_g36249 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_452(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_455(0), ZN => gl_rom_n_168);
  gl_rom_g36250 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_764(1), B1 => FE_OFN19_gl_rom_n_21, B2 => gl_rom_rom_761(1), ZN => gl_rom_n_167);
  gl_rom_g36251 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_450(0), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_454(0), ZN => gl_rom_n_166);
  gl_rom_g36252 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_762(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_767(1), ZN => gl_rom_n_165);
  gl_rom_g36253 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_760(1), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_763(1), ZN => gl_rom_n_164);
  gl_rom_g36254 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_728(0), B1 => FE_OFN6_gl_rom_n_18, B2 => gl_rom_rom_732(0), ZN => gl_rom_n_163);
  gl_rom_g36255 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_449(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_453(0), ZN => gl_rom_n_162);
  gl_rom_g36256 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_746(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_751(1), ZN => gl_rom_n_161);
  gl_rom_g36257 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_748(1), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_750(1), ZN => gl_rom_n_160);
  gl_rom_g36258 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_448(0), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_451(0), ZN => gl_rom_n_159);
  gl_rom_g36259 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_22, A2 => gl_rom_rom_749(1), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_747(1), ZN => gl_rom_n_158);
  gl_rom_g36260 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_744(1), B1 => FE_OFN19_gl_rom_n_21, B2 => gl_rom_rom_745(1), ZN => gl_rom_n_157);
  gl_rom_g36261 : AOI22D0BWP7T port map(A1 => FE_OFN4_gl_rom_n_16, A2 => gl_rom_rom_758(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_757(1), ZN => gl_rom_n_156);
  gl_rom_g36262 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_756(1), B1 => gl_rom_n_21, B2 => gl_rom_rom_753(1), ZN => gl_rom_n_155);
  gl_rom_g36263 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_738(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_743(0), ZN => gl_rom_n_154);
  gl_rom_g36264 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_444(0), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_447(0), ZN => gl_rom_n_153);
  gl_rom_g36265 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_754(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_759(1), ZN => gl_rom_n_152);
  gl_rom_g36266 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_858(0), B1 => FE_OFN17_gl_rom_n_15, B2 => gl_rom_rom_859(0), ZN => gl_rom_n_151);
  gl_rom_g36267 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_752(1), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_755(1), ZN => gl_rom_n_150);
  gl_rom_g36268 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_442(0), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_446(0), ZN => gl_rom_n_149);
  gl_rom_g36269 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_740(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_742(0), ZN => gl_rom_n_148);
  gl_rom_g36270 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_21, A2 => gl_rom_rom_721(1), B1 => FE_OFN11_gl_rom_n_22, B2 => gl_rom_rom_725(1), ZN => gl_rom_n_147);
  gl_rom_g36271 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_724(1), B1 => FE_OFN4_gl_rom_n_16, B2 => gl_rom_rom_726(1), ZN => gl_rom_n_146);
  gl_rom_g36272 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_441(0), B1 => FE_OFN11_gl_rom_n_22, B2 => gl_rom_rom_445(0), ZN => gl_rom_n_145);
  gl_rom_g36273 : AOI22D0BWP7T port map(A1 => gl_rom_n_22, A2 => gl_rom_rom_965(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_963(0), ZN => gl_rom_n_144);
  gl_rom_g36274 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_722(1), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_723(1), ZN => gl_rom_n_143);
  gl_rom_g36275 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_720(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_727(1), ZN => gl_rom_n_142);
  gl_rom_g36276 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_440(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_443(0), ZN => gl_rom_n_141);
  gl_rom_g36277 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_856(0), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_863(0), ZN => gl_rom_n_140);
  gl_rom_g36278 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_22, A2 => gl_rom_rom_741(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_739(0), ZN => gl_rom_n_139);
  gl_rom_g36279 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_730(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_735(1), ZN => gl_rom_n_138);
  gl_rom_g36280 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_732(1), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_734(1), ZN => gl_rom_n_137);
  gl_rom_g36281 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_425(0), B1 => FE_OFN11_gl_rom_n_22, B2 => gl_rom_rom_429(0), ZN => gl_rom_n_136);
  gl_rom_g36282 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_22, A2 => gl_rom_rom_733(1), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_731(1), ZN => gl_rom_n_135);
  gl_rom_g36283 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_428(0), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_430(0), ZN => gl_rom_n_134);
  gl_rom_g36284 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_728(1), B1 => FE_OFN19_gl_rom_n_21, B2 => gl_rom_rom_729(1), ZN => gl_rom_n_133);
  gl_rom_g36285 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_736(0), B1 => FE_OFN19_gl_rom_n_21, B2 => gl_rom_rom_737(0), ZN => gl_rom_n_132);
  gl_rom_g36286 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_738(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_743(1), ZN => gl_rom_n_131);
  gl_rom_g36287 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_426(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_427(0), ZN => gl_rom_n_130);
  gl_rom_g36288 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_740(1), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_742(1), ZN => gl_rom_n_129);
  gl_rom_g36289 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_22, A2 => gl_rom_rom_741(1), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_739(1), ZN => gl_rom_n_128);
  gl_rom_g36290 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_424(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_431(0), ZN => gl_rom_n_127);
  gl_rom_g36291 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_736(1), B1 => FE_OFN19_gl_rom_n_21, B2 => gl_rom_rom_737(1), ZN => gl_rom_n_126);
  gl_rom_g36292 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_714(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_719(1), ZN => gl_rom_n_125);
  gl_rom_g36293 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_716(1), B1 => FE_OFN4_gl_rom_n_16, B2 => gl_rom_rom_718(1), ZN => gl_rom_n_124);
  gl_rom_g36294 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_412(0), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_415(0), ZN => gl_rom_n_123);
  gl_rom_g36295 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_21, A2 => gl_rom_rom_761(0), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_765(0), ZN => gl_rom_n_122);
  gl_rom_g36296 : AOI22D0BWP7T port map(A1 => FE_OFN11_gl_rom_n_22, A2 => gl_rom_rom_717(1), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_715(1), ZN => gl_rom_n_121);
  gl_rom_g36297 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_712(1), B1 => FE_OFN19_gl_rom_n_21, B2 => gl_rom_rom_713(1), ZN => gl_rom_n_120);
  gl_rom_g36298 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_865(0), B1 => FE_OFN11_gl_rom_n_22, B2 => gl_rom_rom_869(0), ZN => gl_rom_n_119);
  gl_rom_g36299 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_410(0), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_414(0), ZN => gl_rom_n_118);
  gl_rom_g36300 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_706(1), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_711(1), ZN => gl_rom_n_117);
  gl_rom_g36301 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_960(0), B1 => gl_rom_n_21, B2 => gl_rom_rom_961(0), ZN => gl_rom_n_116);
  gl_rom_g36302 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_21, A2 => gl_rom_rom_705(1), B1 => FE_OFN11_gl_rom_n_22, B2 => gl_rom_rom_709(1), ZN => gl_rom_n_115);
  gl_rom_g36303 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_764(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_766(0), ZN => gl_rom_n_114);
  gl_rom_g36304 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_409(0), B1 => FE_OFN11_gl_rom_n_22, B2 => gl_rom_rom_413(0), ZN => gl_rom_n_113);
  gl_rom_g36305 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_408(0), B1 => FE_OFN15_gl_rom_n_15, B2 => gl_rom_rom_411(0), ZN => gl_rom_n_112);
  gl_rom_g36306 : AOI22D0BWP7T port map(A1 => FE_OFN1_gl_rom_n_16, A2 => gl_rom_rom_710(1), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_707(1), ZN => gl_rom_n_111);
  gl_rom_g36307 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_704(1), B1 => FE_OFN7_gl_rom_n_18, B2 => gl_rom_rom_708(1), ZN => gl_rom_n_110);
  gl_rom_g36308 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_868(0), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_870(0), ZN => gl_rom_n_109);
  gl_rom_g36309 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_826(1), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_831(1), ZN => gl_rom_n_108);
  gl_rom_g36310 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_762(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_763(0), ZN => gl_rom_n_107);
  gl_rom_g36311 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_420(0), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_423(0), ZN => gl_rom_n_106);
  gl_rom_g36312 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_825(1), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_829(1), ZN => gl_rom_n_105);
  gl_rom_g36313 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_418(0), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_422(0), ZN => gl_rom_n_104);
  gl_rom_g36314 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_828(1), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_830(1), ZN => gl_rom_n_103);
  gl_rom_g36315 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_824(1), B1 => FE_OFN17_gl_rom_n_15, B2 => gl_rom_rom_827(1), ZN => gl_rom_n_102);
  gl_rom_g36316 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_760(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_767(0), ZN => gl_rom_n_101);
  gl_rom_g36317 : AOI22D0BWP7T port map(A1 => FE_OFN1_gl_rom_n_16, A2 => gl_rom_rom_814(1), B1 => FE_OFN13_gl_rom_n_22, B2 => gl_rom_rom_813(1), ZN => gl_rom_n_100);
  gl_rom_g36318 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_417(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_421(0), ZN => gl_rom_n_99);
  gl_rom_g36319 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_812(1), B1 => FE_OFN20_gl_rom_n_21, B2 => gl_rom_rom_809(1), ZN => gl_rom_n_98);
  gl_rom_g36320 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_416(0), B1 => FE_OFN17_gl_rom_n_15, B2 => gl_rom_rom_419(0), ZN => gl_rom_n_97);
  gl_rom_g36321 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_810(1), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_815(1), ZN => gl_rom_n_96);
  gl_rom_g36322 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_808(1), B1 => FE_OFN17_gl_rom_n_15, B2 => gl_rom_rom_811(1), ZN => gl_rom_n_95);
  gl_rom_g36323 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_796(1), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_799(1), ZN => gl_rom_n_94);
  gl_rom_g36324 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_994(0), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_999(0), ZN => gl_rom_n_93);
  gl_rom_g36325 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_794(1), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_798(1), ZN => gl_rom_n_92);
  gl_rom_g36326 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_866(0), B1 => FE_OFN17_gl_rom_n_15, B2 => gl_rom_rom_867(0), ZN => gl_rom_n_91);
  gl_rom_g36327 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_436(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_439(0), ZN => gl_rom_n_90);
  gl_rom_g36328 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_746(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_751(0), ZN => gl_rom_n_89);
  gl_rom_g36329 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_793(1), B1 => FE_OFN11_gl_rom_n_22, B2 => gl_rom_rom_797(1), ZN => gl_rom_n_88);
  gl_rom_g36330 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_792(1), B1 => FE_OFN17_gl_rom_n_15, B2 => gl_rom_rom_795(1), ZN => gl_rom_n_87);
  gl_rom_g36331 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_434(0), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_438(0), ZN => gl_rom_n_86);
  gl_rom_g36332 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_748(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_750(0), ZN => gl_rom_n_85);
  gl_rom_g36333 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_804(1), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_807(1), ZN => gl_rom_n_84);
  gl_rom_g36334 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_802(1), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_806(1), ZN => gl_rom_n_83);
  gl_rom_g36335 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_21, A2 => gl_rom_rom_433(0), B1 => FE_OFN11_gl_rom_n_22, B2 => gl_rom_rom_437(0), ZN => gl_rom_n_82);
  gl_rom_g36336 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_801(1), B1 => FE_OFN11_gl_rom_n_22, B2 => gl_rom_rom_805(1), ZN => gl_rom_n_81);
  gl_rom_g36337 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_800(1), B1 => FE_OFN17_gl_rom_n_15, B2 => gl_rom_rom_803(1), ZN => gl_rom_n_80);
  gl_rom_g36338 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_432(0), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_435(0), ZN => gl_rom_n_79);
  gl_rom_g36339 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_1010(0), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_1015(0), ZN => gl_rom_n_78);
  gl_rom_g36340 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_22, A2 => gl_rom_rom_749(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_747(0), ZN => gl_rom_n_77);
  gl_rom_g36341 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_818(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_823(1), ZN => gl_rom_n_76);
  gl_rom_g36342 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_864(0), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_871(0), ZN => gl_rom_n_75);
  gl_rom_g36343 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_404(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_407(0), ZN => gl_rom_n_74);
  gl_rom_g36344 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_817(1), B1 => FE_OFN11_gl_rom_n_22, B2 => gl_rom_rom_821(1), ZN => gl_rom_n_73);
  gl_rom_g36345 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_996(0), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_998(0), ZN => gl_rom_n_72);
  gl_rom_g36346 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_820(1), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_822(1), ZN => gl_rom_n_71);
  gl_rom_g36347 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_402(0), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_406(0), ZN => gl_rom_n_70);
  gl_rom_g36348 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_816(1), B1 => FE_OFN17_gl_rom_n_15, B2 => gl_rom_rom_819(1), ZN => gl_rom_n_69);
  gl_rom_g36349 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_744(0), B1 => FE_OFN19_gl_rom_n_21, B2 => gl_rom_rom_745(0), ZN => gl_rom_n_68);
  gl_rom_g36350 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_788(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_791(1), ZN => gl_rom_n_67);
  gl_rom_g36351 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_786(1), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_790(1), ZN => gl_rom_n_66);
  gl_rom_g36352 : AOI22D0BWP7T port map(A1 => FE_OFN19_gl_rom_n_21, A2 => gl_rom_rom_401(0), B1 => FE_OFN11_gl_rom_n_22, B2 => gl_rom_rom_405(0), ZN => gl_rom_n_65);
  gl_rom_g36353 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_785(1), B1 => FE_OFN11_gl_rom_n_22, B2 => gl_rom_rom_789(1), ZN => gl_rom_n_64);
  gl_rom_g36354 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_400(0), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_403(0), ZN => gl_rom_n_63);
  gl_rom_g36355 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_784(1), B1 => FE_OFN17_gl_rom_n_15, B2 => gl_rom_rom_787(1), ZN => gl_rom_n_62);
  gl_rom_g36356 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_777(1), B1 => FE_OFN11_gl_rom_n_22, B2 => gl_rom_rom_781(1), ZN => gl_rom_n_61);
  gl_rom_g36357 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_780(1), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_782(1), ZN => gl_rom_n_60);
  gl_rom_g36358 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_396(0), B1 => FE_OFN10_gl_rom_n_17, B2 => gl_rom_rom_399(0), ZN => gl_rom_n_59);
  gl_rom_g36359 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_714(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_719(0), ZN => gl_rom_n_58);
  gl_rom_g36360 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_778(1), B1 => FE_OFN17_gl_rom_n_15, B2 => gl_rom_rom_779(1), ZN => gl_rom_n_57);
  gl_rom_g36361 : AOI22D0BWP7T port map(A1 => FE_OFN29_gl_rom_n_20, A2 => gl_rom_rom_394(0), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_398(0), ZN => gl_rom_n_56);
  gl_rom_g36362 : AOI22D0BWP7T port map(A1 => FE_OFN25_gl_rom_n_19, A2 => gl_rom_rom_776(1), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_783(1), ZN => gl_rom_n_55);
  gl_rom_g36363 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_772(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_775(1), ZN => gl_rom_n_54);
  gl_rom_g36364 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_716(0), B1 => FE_OFN3_gl_rom_n_16, B2 => gl_rom_rom_718(0), ZN => gl_rom_n_53);
  gl_rom_g36365 : AOI22D0BWP7T port map(A1 => gl_rom_n_21, A2 => gl_rom_rom_393(0), B1 => gl_rom_n_22, B2 => gl_rom_rom_397(0), ZN => gl_rom_n_52);
  gl_rom_g36366 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_770(1), B1 => FE_OFN1_gl_rom_n_16, B2 => gl_rom_rom_774(1), ZN => gl_rom_n_51);
  gl_rom_g36367 : AOI22D0BWP7T port map(A1 => FE_OFN1_gl_rom_n_16, A2 => gl_rom_rom_886(0), B1 => FE_OFN11_gl_rom_n_22, B2 => gl_rom_rom_885(0), ZN => gl_rom_n_50);
  gl_rom_g36368 : AOI22D0BWP7T port map(A1 => FE_OFN26_gl_rom_n_19, A2 => gl_rom_rom_392(0), B1 => FE_OFN14_gl_rom_n_15, B2 => gl_rom_rom_395(0), ZN => gl_rom_n_49);
  gl_rom_g36369 : AOI22D0BWP7T port map(A1 => FE_OFN20_gl_rom_n_21, A2 => gl_rom_rom_769(1), B1 => FE_OFN11_gl_rom_n_22, B2 => gl_rom_rom_773(1), ZN => gl_rom_n_48);
  gl_rom_g36370 : AOI22D0BWP7T port map(A1 => FE_OFN24_gl_rom_n_19, A2 => gl_rom_rom_768(1), B1 => FE_OFN17_gl_rom_n_15, B2 => gl_rom_rom_771(1), ZN => gl_rom_n_47);
  gl_rom_g36371 : AOI22D0BWP7T port map(A1 => FE_OFN28_gl_rom_n_20, A2 => gl_rom_rom_954(0), B1 => FE_OFN9_gl_rom_n_17, B2 => gl_rom_rom_959(0), ZN => gl_rom_n_46);
  gl_rom_g36372 : AOI22D0BWP7T port map(A1 => FE_OFN6_gl_rom_n_18, A2 => gl_rom_rom_884(0), B1 => FE_OFN19_gl_rom_n_21, B2 => gl_rom_rom_881(0), ZN => gl_rom_n_45);
  gl_rom_g36373 : AOI22D0BWP7T port map(A1 => FE_OFN13_gl_rom_n_22, A2 => gl_rom_rom_717(0), B1 => FE_OFN18_gl_rom_n_15, B2 => gl_rom_rom_715(0), ZN => gl_rom_n_44);
  gl_rom_g36374 : AOI22D0BWP7T port map(A1 => FE_OFN5_gl_rom_n_18, A2 => gl_rom_rom_1012(1), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_1015(1), ZN => gl_rom_n_43);
  gl_rom_g36375 : AOI22D0BWP7T port map(A1 => FE_OFN7_gl_rom_n_18, A2 => gl_rom_rom_388(0), B1 => FE_OFN8_gl_rom_n_17, B2 => gl_rom_rom_391(0), ZN => gl_rom_n_42);
  gl_rom_g36376 : AOI22D0BWP7T port map(A1 => gl_rom_n_20, A2 => gl_rom_rom_1010(1), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_1014(1), ZN => gl_rom_n_41);
  gl_rom_g36377 : AOI22D0BWP7T port map(A1 => FE_OFN27_gl_rom_n_20, A2 => gl_rom_rom_386(0), B1 => FE_OFN0_gl_rom_n_16, B2 => gl_rom_rom_390(0), ZN => gl_rom_n_40);
  gl_rom_g36378 : AOI22D0BWP7T port map(A1 => FE_OFN22_gl_rom_n_21, A2 => gl_rom_rom_1009(1), B1 => gl_rom_n_22, B2 => gl_rom_rom_1013(1), ZN => gl_rom_n_39);
  gl_rom_g36379 : AN2D1BWP7T port map(A1 => gl_rom_n_13, A2 => gl_sig_e(8), Z => gl_rom_n_38);
  gl_rom_g36380 : INR2D1BWP7T port map(A1 => gl_sig_e(8), B1 => gl_rom_n_1, ZN => gl_rom_n_37);
  gl_rom_g36381 : INR2D1BWP7T port map(A1 => gl_sig_e(8), B1 => gl_rom_n_2, ZN => gl_rom_n_36);
  gl_rom_g36382 : NR2D1BWP7T port map(A1 => gl_rom_n_1, A2 => gl_sig_e(8), ZN => gl_rom_n_35);
  gl_rom_g36383 : NR2D1BWP7T port map(A1 => gl_rom_n_9, A2 => gl_sig_e(8), ZN => gl_rom_n_34);
  gl_rom_g36384 : NR2D1BWP7T port map(A1 => gl_rom_n_2, A2 => gl_sig_e(8), ZN => gl_rom_n_33);
  gl_rom_g36385 : INR2D1BWP7T port map(A1 => gl_rom_n_13, B1 => gl_sig_e(8), ZN => gl_rom_n_32);
  gl_rom_g36386 : INR2D1BWP7T port map(A1 => gl_sig_e(8), B1 => gl_rom_n_9, ZN => gl_rom_n_31);
  gl_rom_g36387 : AN2D1BWP7T port map(A1 => gl_rom_n_8, A2 => gl_sig_e(4), Z => gl_rom_n_30);
  gl_rom_g36388 : NR2XD1BWP7T port map(A1 => gl_rom_n_7, A2 => gl_sig_e(4), ZN => gl_rom_n_29);
  gl_rom_g36389 : AN2D1BWP7T port map(A1 => gl_rom_n_4, A2 => gl_sig_e(4), Z => gl_rom_n_28);
  gl_rom_g36390 : INR2D2BWP7T port map(A1 => gl_sig_e(4), B1 => gl_rom_n_11, ZN => gl_rom_n_27);
  gl_rom_g36391 : NR2XD1BWP7T port map(A1 => gl_rom_n_11, A2 => gl_sig_e(4), ZN => gl_rom_n_26);
  gl_rom_g36392 : AN2D1BWP7T port map(A1 => gl_rom_n_14, A2 => gl_sig_e(4), Z => gl_rom_n_25);
  gl_rom_g36393 : INR2D2BWP7T port map(A1 => gl_rom_n_14, B1 => gl_sig_e(4), ZN => gl_rom_n_24);
  gl_rom_g36394 : NR2XD1BWP7T port map(A1 => gl_rom_n_5, A2 => gl_sig_e(4), ZN => gl_rom_n_23);
  gl_rom_g36395 : AN2D2BWP7T port map(A1 => gl_rom_n_3, A2 => gl_sig_e(2), Z => gl_rom_n_22);
  gl_rom_g36396 : AN2D2BWP7T port map(A1 => gl_rom_n_3, A2 => gl_rom_n_0, Z => gl_rom_n_21);
  gl_rom_g36397 : AN2D2BWP7T port map(A1 => gl_rom_n_10, A2 => gl_rom_n_0, Z => gl_rom_n_20);
  gl_rom_g36398 : AN2D2BWP7T port map(A1 => gl_rom_n_6, A2 => gl_rom_n_0, Z => gl_rom_n_19);
  gl_rom_g36399 : AN2D1BWP7T port map(A1 => gl_rom_n_6, A2 => gl_sig_e(2), Z => gl_rom_n_18);
  gl_rom_g36400 : AN2D1BWP7T port map(A1 => gl_rom_n_12, A2 => gl_sig_e(2), Z => gl_rom_n_17);
  gl_rom_g36401 : AN2D1BWP7T port map(A1 => gl_rom_n_10, A2 => gl_sig_e(2), Z => gl_rom_n_16);
  gl_rom_g36402 : AN2D2BWP7T port map(A1 => gl_rom_n_12, A2 => gl_rom_n_0, Z => gl_rom_n_15);
  gl_rom_g36403 : NR2XD0BWP7T port map(A1 => gl_sig_e(5), A2 => gl_sig_e(3), ZN => gl_rom_n_14);
  gl_rom_g36404 : NR2D0BWP7T port map(A1 => gl_sig_e(7), A2 => gl_sig_e(6), ZN => gl_rom_n_13);
  gl_rom_g36405 : AN2D1BWP7T port map(A1 => gl_sig_e(0), A2 => gl_sig_e(1), Z => gl_rom_n_12);
  gl_rom_g36406 : ND2D1BWP7T port map(A1 => gl_sig_e(3), A2 => gl_sig_e(5), ZN => gl_rom_n_11);
  gl_rom_g36407 : INR2D1BWP7T port map(A1 => gl_sig_e(1), B1 => gl_sig_e(0), ZN => gl_rom_n_10);
  gl_rom_g36408 : CKND2D1BWP7T port map(A1 => gl_sig_e(7), A2 => gl_sig_e(6), ZN => gl_rom_n_9);
  gl_rom_g36409 : INVD0BWP7T port map(I => gl_rom_n_7, ZN => gl_rom_n_8);
  gl_rom_g36410 : INVD0BWP7T port map(I => gl_rom_n_4, ZN => gl_rom_n_5);
  gl_rom_g36411 : IND2D1BWP7T port map(A1 => gl_sig_e(5), B1 => gl_sig_e(3), ZN => gl_rom_n_7);
  gl_rom_g36412 : NR2D1BWP7T port map(A1 => gl_sig_e(0), A2 => gl_sig_e(1), ZN => gl_rom_n_6);
  gl_rom_g36413 : INR2D1BWP7T port map(A1 => gl_sig_e(5), B1 => gl_sig_e(3), ZN => gl_rom_n_4);
  gl_rom_g36414 : INR2D1BWP7T port map(A1 => gl_sig_e(0), B1 => gl_sig_e(1), ZN => gl_rom_n_3);
  gl_rom_g36415 : IND2D1BWP7T port map(A1 => gl_sig_e(7), B1 => gl_sig_e(6), ZN => gl_rom_n_2);
  gl_rom_g36416 : IND2D1BWP7T port map(A1 => gl_sig_e(6), B1 => gl_sig_e(7), ZN => gl_rom_n_1);
  gl_rom_g36417 : INVD1BWP7T port map(I => gl_sig_e(2), ZN => gl_rom_n_0);
  gl_ram_g13776 : MOAI22D0BWP7T port map(A1 => gl_ram_n_826, A2 => gl_ram_n_794, B1 => gl_ram_n_822, B2 => gl_ram_n_794, ZN => gl_sig_ram(2));
  gl_ram_g13777 : MOAI22D0BWP7T port map(A1 => gl_ram_n_825, A2 => gl_ram_n_794, B1 => gl_ram_n_821, B2 => gl_ram_n_794, ZN => gl_sig_ram(0));
  gl_ram_g13778 : MOAI22D0BWP7T port map(A1 => gl_ram_n_824, A2 => gl_ram_n_794, B1 => gl_ram_n_823, B2 => gl_ram_n_794, ZN => gl_sig_ram(1));
  gl_ram_g13779 : AN4D0BWP7T port map(A1 => gl_ram_n_819, A2 => gl_ram_n_820, A3 => gl_ram_n_800, A4 => gl_ram_n_810, Z => gl_ram_n_826);
  gl_ram_g13780 : AN4D0BWP7T port map(A1 => gl_ram_n_818, A2 => gl_ram_n_817, A3 => gl_ram_n_799, A4 => gl_ram_n_807, Z => gl_ram_n_825);
  gl_ram_g13781 : AN4D1BWP7T port map(A1 => gl_ram_n_815, A2 => gl_ram_n_816, A3 => gl_ram_n_804, A4 => gl_ram_n_798, Z => gl_ram_n_824);
  gl_ram_g13782 : ND4D0BWP7T port map(A1 => gl_ram_n_802, A2 => gl_ram_n_809, A3 => gl_ram_n_806, A4 => gl_ram_n_811, ZN => gl_ram_n_823);
  gl_ram_g13783 : ND4D0BWP7T port map(A1 => gl_ram_n_801, A2 => gl_ram_n_808, A3 => gl_ram_n_812, A4 => gl_ram_n_814, ZN => gl_ram_n_822);
  gl_ram_g13784 : ND4D0BWP7T port map(A1 => gl_ram_n_805, A2 => gl_ram_n_803, A3 => gl_ram_n_813, A4 => gl_ram_n_797, ZN => gl_ram_n_821);
  gl_ram_g13785 : AOI22D0BWP7T port map(A1 => gl_ram_n_795, A2 => gl_ram_ram_96(2), B1 => gl_ram_n_570, B2 => gl_ram_ram_97(2), ZN => gl_ram_n_820);
  gl_ram_g13786 : AOI22D0BWP7T port map(A1 => gl_ram_n_796, A2 => gl_ram_ram_98(2), B1 => gl_ram_n_569, B2 => gl_ram_ram_99(2), ZN => gl_ram_n_819);
  gl_ram_g13787 : AOI22D0BWP7T port map(A1 => gl_ram_n_796, A2 => gl_ram_ram_98(0), B1 => gl_ram_n_569, B2 => gl_ram_ram_99(0), ZN => gl_ram_n_818);
  gl_ram_g13788 : AOI22D0BWP7T port map(A1 => gl_ram_n_795, A2 => gl_ram_ram_96(0), B1 => gl_ram_n_570, B2 => gl_ram_ram_97(0), ZN => gl_ram_n_817);
  gl_ram_g13789 : AOI22D0BWP7T port map(A1 => gl_ram_n_795, A2 => gl_ram_ram_96(1), B1 => gl_ram_n_570, B2 => gl_ram_ram_97(1), ZN => gl_ram_n_816);
  gl_ram_g13790 : AOI22D0BWP7T port map(A1 => gl_ram_n_796, A2 => gl_ram_ram_98(1), B1 => gl_ram_n_569, B2 => gl_ram_ram_99(1), ZN => gl_ram_n_815);
  gl_ram_g13791 : AOI22D0BWP7T port map(A1 => gl_ram_n_787, A2 => gl_ram_n_749, B1 => gl_ram_n_793, B2 => gl_ram_n_756, ZN => gl_ram_n_814);
  gl_ram_g13792 : AOI22D0BWP7T port map(A1 => gl_ram_n_789, A2 => gl_ram_n_757, B1 => gl_ram_n_788, B2 => gl_ram_n_750, ZN => gl_ram_n_813);
  gl_ram_g13793 : AOI22D0BWP7T port map(A1 => gl_ram_n_789, A2 => gl_ram_n_773, B1 => gl_ram_n_788, B2 => gl_ram_n_741, ZN => gl_ram_n_812);
  gl_ram_g13794 : AOI22D0BWP7T port map(A1 => gl_ram_n_787, A2 => gl_ram_n_774, B1 => gl_ram_n_793, B2 => gl_ram_n_766, ZN => gl_ram_n_811);
  gl_ram_g13795 : AOI22D0BWP7T port map(A1 => gl_ram_n_791, A2 => gl_ram_n_764, B1 => gl_ram_n_785, B2 => gl_ram_n_771, ZN => gl_ram_n_810);
  gl_ram_g13796 : AOI22D0BWP7T port map(A1 => gl_ram_n_791, A2 => gl_ram_n_763, B1 => gl_ram_n_785, B2 => gl_ram_n_765, ZN => gl_ram_n_809);
  gl_ram_g13797 : AOI22D0BWP7T port map(A1 => gl_ram_n_791, A2 => gl_ram_n_759, B1 => gl_ram_n_785, B2 => gl_ram_n_761, ZN => gl_ram_n_808);
  gl_ram_g13798 : AOI22D0BWP7T port map(A1 => gl_ram_n_791, A2 => gl_ram_n_755, B1 => gl_ram_n_785, B2 => gl_ram_n_748, ZN => gl_ram_n_807);
  gl_ram_g13799 : AOI22D0BWP7T port map(A1 => gl_ram_n_789, A2 => gl_ram_n_767, B1 => gl_ram_n_788, B2 => gl_ram_n_768, ZN => gl_ram_n_806);
  gl_ram_g13800 : AOI22D0BWP7T port map(A1 => gl_ram_n_786, A2 => gl_ram_n_744, B1 => gl_ram_n_792, B2 => gl_ram_n_746, ZN => gl_ram_n_805);
  gl_ram_g13801 : AOI22D0BWP7T port map(A1 => gl_ram_n_791, A2 => gl_ram_n_743, B1 => gl_ram_n_785, B2 => gl_ram_n_747, ZN => gl_ram_n_804);
  gl_ram_g13802 : AOI22D0BWP7T port map(A1 => gl_ram_n_791, A2 => gl_ram_n_740, B1 => gl_ram_n_785, B2 => gl_ram_n_742, ZN => gl_ram_n_803);
  gl_ram_g13803 : AOI22D0BWP7T port map(A1 => gl_ram_n_786, A2 => gl_ram_n_770, B1 => gl_ram_n_792, B2 => gl_ram_n_772, ZN => gl_ram_n_802);
  gl_ram_g13804 : AOI22D0BWP7T port map(A1 => gl_ram_n_786, A2 => gl_ram_n_775, B1 => gl_ram_n_792, B2 => gl_ram_n_769, ZN => gl_ram_n_801);
  gl_ram_g13805 : AOI22D0BWP7T port map(A1 => gl_ram_n_786, A2 => gl_ram_n_745, B1 => gl_ram_n_792, B2 => gl_ram_n_762, ZN => gl_ram_n_800);
  gl_ram_g13806 : AOI22D0BWP7T port map(A1 => gl_ram_n_786, A2 => gl_ram_n_758, B1 => gl_ram_n_792, B2 => gl_ram_n_760, ZN => gl_ram_n_799);
  gl_ram_g13807 : AOI22D0BWP7T port map(A1 => gl_ram_n_786, A2 => gl_ram_n_751, B1 => gl_ram_n_792, B2 => gl_ram_n_754, ZN => gl_ram_n_798);
  gl_ram_g13808 : AOI22D0BWP7T port map(A1 => gl_ram_n_787, A2 => gl_ram_n_752, B1 => gl_ram_n_793, B2 => gl_ram_n_753, ZN => gl_ram_n_797);
  gl_ram_g13809 : NR2D0BWP7T port map(A1 => gl_ram_n_790, A2 => gl_ram_n_591, ZN => gl_ram_n_796);
  gl_ram_g13810 : NR2D0BWP7T port map(A1 => gl_ram_n_790, A2 => gl_ram_n_589, ZN => gl_ram_n_795);
  gl_ram_g13813 : XNR2D1BWP7T port map(A1 => gl_ram_n_782, A2 => gl_sig_y(3), ZN => gl_ram_n_794);
  gl_ram_g13814 : INVD0BWP7T port map(I => gl_ram_n_790, ZN => gl_ram_n_789);
  gl_ram_g13815 : NR2D0BWP7T port map(A1 => gl_ram_n_783, A2 => gl_ram_n_778, ZN => gl_ram_n_793);
  gl_ram_g13816 : NR2D0BWP7T port map(A1 => gl_ram_n_784, A2 => gl_ram_n_778, ZN => gl_ram_n_792);
  gl_ram_g13817 : INR2D0BWP7T port map(A1 => gl_ram_n_779, B1 => gl_ram_n_784, ZN => gl_ram_n_791);
  gl_ram_g13818 : ND2D0BWP7T port map(A1 => gl_ram_n_784, A2 => gl_ram_n_779, ZN => gl_ram_n_790);
  gl_ram_g13819 : NR2D0BWP7T port map(A1 => gl_ram_n_783, A2 => gl_ram_n_781, ZN => gl_ram_n_788);
  gl_ram_g13820 : NR2D0BWP7T port map(A1 => gl_ram_n_783, A2 => gl_ram_n_780, ZN => gl_ram_n_787);
  gl_ram_g13821 : NR2D0BWP7T port map(A1 => gl_ram_n_784, A2 => gl_ram_n_781, ZN => gl_ram_n_786);
  gl_ram_g13822 : NR2D0BWP7T port map(A1 => gl_ram_n_784, A2 => gl_ram_n_780, ZN => gl_ram_n_785);
  gl_ram_g13823 : CKND1BWP7T port map(I => gl_ram_n_784, ZN => gl_ram_n_783);
  gl_ram_g13824 : FA1D0BWP7T port map(A => gl_ram_n_573, B => gl_sig_y(2), CI => gl_ram_n_776, CO => gl_ram_n_782, S => gl_ram_n_784);
  gl_ram_g13825 : IND2D0BWP7T port map(A1 => gl_ram_n_777, B1 => gl_ram_n_739, ZN => gl_ram_n_781);
  gl_ram_g13826 : IND2D0BWP7T port map(A1 => gl_ram_n_739, B1 => gl_ram_n_777, ZN => gl_ram_n_780);
  gl_ram_g13827 : NR2D0BWP7T port map(A1 => gl_ram_n_777, A2 => gl_ram_n_739, ZN => gl_ram_n_779);
  gl_ram_g13828 : ND2D0BWP7T port map(A1 => gl_ram_n_777, A2 => gl_ram_n_739, ZN => gl_ram_n_778);
  gl_ram_g13829 : FA1D0BWP7T port map(A => gl_ram_n_574, B => gl_ram_n_575, CI => gl_ram_n_738, CO => gl_ram_n_776, S => gl_ram_n_777);
  gl_ram_g13830 : ND4D0BWP7T port map(A1 => gl_ram_n_693, A2 => gl_ram_n_684, A3 => gl_ram_n_695, A4 => gl_ram_n_689, ZN => gl_ram_n_775);
  gl_ram_g13831 : ND4D0BWP7T port map(A1 => gl_ram_n_727, A2 => gl_ram_n_724, A3 => gl_ram_n_728, A4 => gl_ram_n_726, ZN => gl_ram_n_774);
  gl_ram_g13832 : ND4D0BWP7T port map(A1 => gl_ram_n_723, A2 => gl_ram_n_716, A3 => gl_ram_n_725, A4 => gl_ram_n_720, ZN => gl_ram_n_773);
  gl_ram_g13833 : ND4D0BWP7T port map(A1 => gl_ram_n_721, A2 => gl_ram_n_717, A3 => gl_ram_n_722, A4 => gl_ram_n_719, ZN => gl_ram_n_772);
  gl_ram_g13834 : ND4D0BWP7T port map(A1 => gl_ram_n_711, A2 => gl_ram_n_698, A3 => gl_ram_n_718, A4 => gl_ram_n_705, ZN => gl_ram_n_771);
  gl_ram_g13835 : ND4D0BWP7T port map(A1 => gl_ram_n_712, A2 => gl_ram_n_709, A3 => gl_ram_n_715, A4 => gl_ram_n_714, ZN => gl_ram_n_770);
  gl_ram_g13836 : ND4D0BWP7T port map(A1 => gl_ram_n_704, A2 => gl_ram_n_700, A3 => gl_ram_n_710, A4 => gl_ram_n_708, ZN => gl_ram_n_769);
  gl_ram_g13837 : ND4D0BWP7T port map(A1 => gl_ram_n_703, A2 => gl_ram_n_702, A3 => gl_ram_n_707, A4 => gl_ram_n_706, ZN => gl_ram_n_768);
  gl_ram_g13838 : ND4D0BWP7T port map(A1 => gl_ram_n_697, A2 => gl_ram_n_694, A3 => gl_ram_n_699, A4 => gl_ram_n_696, ZN => gl_ram_n_767);
  gl_ram_g13839 : ND4D0BWP7T port map(A1 => gl_ram_n_732, A2 => gl_ram_n_730, A3 => gl_ram_n_735, A4 => gl_ram_n_734, ZN => gl_ram_n_766);
  gl_ram_g13840 : ND4D0BWP7T port map(A1 => gl_ram_n_690, A2 => gl_ram_n_686, A3 => gl_ram_n_692, A4 => gl_ram_n_688, ZN => gl_ram_n_765);
  gl_ram_g13841 : ND4D0BWP7T port map(A1 => gl_ram_n_675, A2 => gl_ram_n_668, A3 => gl_ram_n_685, A4 => gl_ram_n_673, ZN => gl_ram_n_764);
  gl_ram_g13842 : ND4D0BWP7T port map(A1 => gl_ram_n_681, A2 => gl_ram_n_677, A3 => gl_ram_n_682, A4 => gl_ram_n_680, ZN => gl_ram_n_763);
  gl_ram_g13843 : ND4D0BWP7T port map(A1 => gl_ram_n_737, A2 => gl_ram_n_632, A3 => gl_ram_n_676, A4 => gl_ram_n_651, ZN => gl_ram_n_762);
  gl_ram_g13844 : ND4D0BWP7T port map(A1 => gl_ram_n_674, A2 => gl_ram_n_671, A3 => gl_ram_n_679, A4 => gl_ram_n_678, ZN => gl_ram_n_761);
  gl_ram_g13845 : ND4D0BWP7T port map(A1 => gl_ram_n_669, A2 => gl_ram_n_667, A3 => gl_ram_n_672, A4 => gl_ram_n_670, ZN => gl_ram_n_760);
  gl_ram_g13846 : ND4D0BWP7T port map(A1 => gl_ram_n_662, A2 => gl_ram_n_657, A3 => gl_ram_n_594, A4 => gl_ram_n_659, ZN => gl_ram_n_759);
  gl_ram_g13847 : ND4D0BWP7T port map(A1 => gl_ram_n_663, A2 => gl_ram_n_660, A3 => gl_ram_n_664, A4 => gl_ram_n_661, ZN => gl_ram_n_758);
  gl_ram_g13848 : ND4D0BWP7T port map(A1 => gl_ram_n_621, A2 => gl_ram_n_619, A3 => gl_ram_n_623, A4 => gl_ram_n_620, ZN => gl_ram_n_757);
  gl_ram_g13849 : ND4D0BWP7T port map(A1 => gl_ram_n_647, A2 => gl_ram_n_635, A3 => gl_ram_n_653, A4 => gl_ram_n_643, ZN => gl_ram_n_756);
  gl_ram_g13850 : ND4D0BWP7T port map(A1 => gl_ram_n_650, A2 => gl_ram_n_648, A3 => gl_ram_n_652, A4 => gl_ram_n_649, ZN => gl_ram_n_755);
  gl_ram_g13851 : ND4D0BWP7T port map(A1 => gl_ram_n_642, A2 => gl_ram_n_636, A3 => gl_ram_n_645, A4 => gl_ram_n_639, ZN => gl_ram_n_754);
  gl_ram_g13852 : ND4D0BWP7T port map(A1 => gl_ram_n_641, A2 => gl_ram_n_640, A3 => gl_ram_n_646, A4 => gl_ram_n_644, ZN => gl_ram_n_753);
  gl_ram_g13853 : ND4D0BWP7T port map(A1 => gl_ram_n_637, A2 => gl_ram_n_633, A3 => gl_ram_n_638, A4 => gl_ram_n_634, ZN => gl_ram_n_752);
  gl_ram_g13854 : ND4D0BWP7T port map(A1 => gl_ram_n_628, A2 => gl_ram_n_622, A3 => gl_ram_n_630, A4 => gl_ram_n_624, ZN => gl_ram_n_751);
  gl_ram_g13855 : ND4D0BWP7T port map(A1 => gl_ram_n_629, A2 => gl_ram_n_626, A3 => gl_ram_n_631, A4 => gl_ram_n_627, ZN => gl_ram_n_750);
  gl_ram_g13856 : ND4D0BWP7T port map(A1 => gl_ram_n_618, A2 => gl_ram_n_687, A3 => gl_ram_n_625, A4 => gl_ram_n_612, ZN => gl_ram_n_749);
  gl_ram_g13857 : ND4D0BWP7T port map(A1 => gl_ram_n_656, A2 => gl_ram_n_654, A3 => gl_ram_n_658, A4 => gl_ram_n_655, ZN => gl_ram_n_748);
  gl_ram_g13858 : ND4D0BWP7T port map(A1 => gl_ram_n_614, A2 => gl_ram_n_609, A3 => gl_ram_n_617, A4 => gl_ram_n_691, ZN => gl_ram_n_747);
  gl_ram_g13859 : ND4D0BWP7T port map(A1 => gl_ram_n_683, A2 => gl_ram_n_613, A3 => gl_ram_n_616, A4 => gl_ram_n_615, ZN => gl_ram_n_746);
  gl_ram_g13860 : ND4D0BWP7T port map(A1 => gl_ram_n_666, A2 => gl_ram_n_729, A3 => gl_ram_n_701, A4 => gl_ram_n_603, ZN => gl_ram_n_745);
  gl_ram_g13861 : ND4D0BWP7T port map(A1 => gl_ram_n_610, A2 => gl_ram_n_607, A3 => gl_ram_n_611, A4 => gl_ram_n_608, ZN => gl_ram_n_744);
  gl_ram_g13862 : ND4D0BWP7T port map(A1 => gl_ram_n_713, A2 => gl_ram_n_665, A3 => gl_ram_n_606, A4 => gl_ram_n_602, ZN => gl_ram_n_743);
  gl_ram_g13863 : ND4D0BWP7T port map(A1 => gl_ram_n_601, A2 => gl_ram_n_600, A3 => gl_ram_n_605, A4 => gl_ram_n_604, ZN => gl_ram_n_742);
  gl_ram_g13864 : ND4D0BWP7T port map(A1 => gl_ram_n_736, A2 => gl_ram_n_731, A3 => gl_ram_n_598, A4 => gl_ram_n_733, ZN => gl_ram_n_741);
  gl_ram_g13865 : ND4D0BWP7T port map(A1 => gl_ram_n_597, A2 => gl_ram_n_595, A3 => gl_ram_n_599, A4 => gl_ram_n_596, ZN => gl_ram_n_740);
  gl_ram_g13866 : FA1D0BWP7T port map(A => gl_ram_n_576, B => gl_sig_y(2), CI => gl_ram_n_581, CO => gl_ram_n_738, S => gl_ram_n_739);
  gl_ram_g13867 : AOI22D0BWP7T port map(A1 => gl_ram_ram_88(2), A2 => gl_ram_n_590, B1 => gl_ram_ram_91(2), B2 => gl_ram_n_584, ZN => gl_ram_n_737);
  gl_ram_g13868 : AOI22D0BWP7T port map(A1 => gl_ram_ram_41(2), A2 => gl_ram_n_588, B1 => gl_ram_ram_42(2), B2 => gl_ram_n_592, ZN => gl_ram_n_736);
  gl_ram_g13869 : AOI22D0BWP7T port map(A1 => gl_ram_ram_62(1), A2 => gl_ram_n_593, B1 => gl_ram_ram_63(1), B2 => gl_ram_n_587, ZN => gl_ram_n_735);
  gl_ram_g13870 : AOI22D0BWP7T port map(A1 => gl_ram_ram_60(1), A2 => gl_ram_n_586, B1 => gl_ram_ram_61(1), B2 => gl_ram_n_585, ZN => gl_ram_n_734);
  gl_ram_g13871 : AOI22D0BWP7T port map(A1 => gl_ram_ram_44(2), A2 => gl_ram_n_586, B1 => gl_ram_ram_45(2), B2 => gl_ram_n_585, ZN => gl_ram_n_733);
  gl_ram_g13872 : AOI22D0BWP7T port map(A1 => gl_ram_ram_57(1), A2 => gl_ram_n_588, B1 => gl_ram_ram_58(1), B2 => gl_ram_n_592, ZN => gl_ram_n_732);
  gl_ram_g13873 : AOI22D0BWP7T port map(A1 => gl_ram_ram_40(2), A2 => gl_ram_n_590, B1 => FE_PHN512_gl_ram_ram_43_2, B2 => gl_ram_n_584, ZN => gl_ram_n_731);
  gl_ram_g13874 : AOI22D0BWP7T port map(A1 => gl_ram_ram_56(1), A2 => gl_ram_n_590, B1 => gl_ram_ram_59(1), B2 => gl_ram_n_584, ZN => gl_ram_n_730);
  gl_ram_g13875 : AOI22D0BWP7T port map(A1 => gl_ram_ram_72(2), A2 => gl_ram_n_590, B1 => gl_ram_ram_75(2), B2 => gl_ram_n_584, ZN => gl_ram_n_729);
  gl_ram_g13876 : AOI22D0BWP7T port map(A1 => gl_ram_ram_54(1), A2 => gl_ram_n_593, B1 => gl_ram_ram_55(1), B2 => gl_ram_n_587, ZN => gl_ram_n_728);
  gl_ram_g13877 : AOI22D0BWP7T port map(A1 => gl_ram_ram_49(1), A2 => gl_ram_n_588, B1 => gl_ram_ram_50(1), B2 => gl_ram_n_592, ZN => gl_ram_n_727);
  gl_ram_g13878 : AOI22D0BWP7T port map(A1 => gl_ram_ram_52(1), A2 => gl_ram_n_586, B1 => gl_ram_ram_53(1), B2 => gl_ram_n_585, ZN => gl_ram_n_726);
  gl_ram_g13879 : AOI22D0BWP7T port map(A1 => gl_ram_ram_38(2), A2 => gl_ram_n_593, B1 => gl_ram_ram_39(2), B2 => gl_ram_n_587, ZN => gl_ram_n_725);
  gl_ram_g13880 : AOI22D0BWP7T port map(A1 => gl_ram_ram_48(1), A2 => gl_ram_n_590, B1 => gl_ram_ram_51(1), B2 => gl_ram_n_584, ZN => gl_ram_n_724);
  gl_ram_g13881 : AOI22D0BWP7T port map(A1 => gl_ram_ram_33(2), A2 => gl_ram_n_588, B1 => gl_ram_ram_34(2), B2 => gl_ram_n_592, ZN => gl_ram_n_723);
  gl_ram_g13882 : AOI22D0BWP7T port map(A1 => gl_ram_ram_30(1), A2 => gl_ram_n_593, B1 => gl_ram_ram_31(1), B2 => gl_ram_n_587, ZN => gl_ram_n_722);
  gl_ram_g13883 : AOI22D0BWP7T port map(A1 => gl_ram_ram_24(1), A2 => gl_ram_n_590, B1 => gl_ram_ram_27(1), B2 => gl_ram_n_584, ZN => gl_ram_n_721);
  gl_ram_g13884 : AOI22D0BWP7T port map(A1 => gl_ram_ram_36(2), A2 => gl_ram_n_586, B1 => gl_ram_ram_37(2), B2 => gl_ram_n_585, ZN => gl_ram_n_720);
  gl_ram_g13885 : AOI22D0BWP7T port map(A1 => gl_ram_ram_28(1), A2 => gl_ram_n_586, B1 => gl_ram_ram_29(1), B2 => gl_ram_n_585, ZN => gl_ram_n_719);
  gl_ram_g13886 : AOI22D0BWP7T port map(A1 => gl_ram_ram_86(2), A2 => gl_ram_n_593, B1 => gl_ram_ram_87(2), B2 => gl_ram_n_587, ZN => gl_ram_n_718);
  gl_ram_g13887 : AOI22D0BWP7T port map(A1 => gl_ram_ram_25(1), A2 => gl_ram_n_588, B1 => gl_ram_ram_26(1), B2 => gl_ram_n_592, ZN => gl_ram_n_717);
  gl_ram_g13888 : AOI22D0BWP7T port map(A1 => gl_ram_ram_32(2), A2 => gl_ram_n_590, B1 => gl_ram_ram_35(2), B2 => gl_ram_n_584, ZN => gl_ram_n_716);
  gl_ram_g13889 : AOI22D0BWP7T port map(A1 => gl_ram_ram_14(1), A2 => gl_ram_n_593, B1 => gl_ram_ram_15(1), B2 => gl_ram_n_587, ZN => gl_ram_n_715);
  gl_ram_g13890 : AOI22D0BWP7T port map(A1 => gl_ram_ram_12(1), A2 => gl_ram_n_586, B1 => gl_ram_ram_13(1), B2 => gl_ram_n_585, ZN => gl_ram_n_714);
  gl_ram_g13891 : AOI22D0BWP7T port map(A1 => gl_ram_ram_66(1), A2 => gl_ram_n_592, B1 => gl_ram_ram_67(1), B2 => gl_ram_n_584, ZN => gl_ram_n_713);
  gl_ram_g13892 : AOI22D0BWP7T port map(A1 => gl_ram_ram_10(1), A2 => gl_ram_n_592, B1 => gl_ram_ram_11(1), B2 => gl_ram_n_584, ZN => gl_ram_n_712);
  gl_ram_g13893 : AOI22D0BWP7T port map(A1 => gl_ram_ram_80(2), A2 => gl_ram_n_590, B1 => gl_ram_ram_83(2), B2 => gl_ram_n_584, ZN => gl_ram_n_711);
  gl_ram_g13894 : AOI22D0BWP7T port map(A1 => gl_ram_ram_30(2), A2 => gl_ram_n_593, B1 => gl_ram_ram_31(2), B2 => gl_ram_n_587, ZN => gl_ram_n_710);
  gl_ram_g13895 : AOI22D0BWP7T port map(A1 => gl_ram_ram_8(1), A2 => gl_ram_n_590, B1 => gl_ram_ram_9(1), B2 => gl_ram_n_588, ZN => gl_ram_n_709);
  gl_ram_g13896 : AOI22D0BWP7T port map(A1 => gl_ram_ram_28(2), A2 => gl_ram_n_586, B1 => gl_ram_ram_29(2), B2 => gl_ram_n_585, ZN => gl_ram_n_708);
  gl_ram_g13897 : AOI22D0BWP7T port map(A1 => gl_ram_ram_46(1), A2 => gl_ram_n_593, B1 => gl_ram_ram_47(1), B2 => gl_ram_n_587, ZN => gl_ram_n_707);
  gl_ram_g13898 : AOI22D0BWP7T port map(A1 => gl_ram_ram_44(1), A2 => gl_ram_n_586, B1 => gl_ram_ram_45(1), B2 => gl_ram_n_585, ZN => gl_ram_n_706);
  gl_ram_g13899 : AOI22D0BWP7T port map(A1 => gl_ram_ram_84(2), A2 => gl_ram_n_586, B1 => gl_ram_ram_85(2), B2 => gl_ram_n_585, ZN => gl_ram_n_705);
  gl_ram_g13900 : AOI22D0BWP7T port map(A1 => gl_ram_ram_25(2), A2 => gl_ram_n_588, B1 => gl_ram_ram_26(2), B2 => gl_ram_n_592, ZN => gl_ram_n_704);
  gl_ram_g13901 : AOI22D0BWP7T port map(A1 => gl_ram_ram_41(1), A2 => gl_ram_n_588, B1 => gl_ram_ram_42(1), B2 => gl_ram_n_592, ZN => gl_ram_n_703);
  gl_ram_g13902 : AOI22D0BWP7T port map(A1 => gl_ram_ram_40(1), A2 => gl_ram_n_590, B1 => FE_PHN658_gl_ram_ram_43_1, B2 => gl_ram_n_584, ZN => gl_ram_n_702);
  gl_ram_g13903 : AOI22D0BWP7T port map(A1 => gl_ram_ram_78(2), A2 => gl_ram_n_593, B1 => gl_ram_ram_79(2), B2 => gl_ram_n_587, ZN => gl_ram_n_701);
  gl_ram_g13904 : AOI22D0BWP7T port map(A1 => gl_ram_ram_24(2), A2 => gl_ram_n_590, B1 => gl_ram_ram_27(2), B2 => gl_ram_n_584, ZN => gl_ram_n_700);
  gl_ram_g13905 : AOI22D0BWP7T port map(A1 => gl_ram_ram_38(1), A2 => gl_ram_n_593, B1 => gl_ram_ram_39(1), B2 => gl_ram_n_587, ZN => gl_ram_n_699);
  gl_ram_g13906 : AOI22D0BWP7T port map(A1 => gl_ram_ram_81(2), A2 => gl_ram_n_588, B1 => gl_ram_ram_82(2), B2 => gl_ram_n_592, ZN => gl_ram_n_698);
  gl_ram_g13907 : AOI22D0BWP7T port map(A1 => gl_ram_ram_33(1), A2 => gl_ram_n_588, B1 => FE_PHN649_gl_ram_ram_34_1, B2 => gl_ram_n_592, ZN => gl_ram_n_697);
  gl_ram_g13908 : AOI22D0BWP7T port map(A1 => gl_ram_ram_36(1), A2 => gl_ram_n_586, B1 => gl_ram_ram_37(1), B2 => gl_ram_n_585, ZN => gl_ram_n_696);
  gl_ram_g13909 : AOI22D0BWP7T port map(A1 => gl_ram_ram_14(2), A2 => gl_ram_n_593, B1 => gl_ram_ram_15(2), B2 => gl_ram_n_587, ZN => gl_ram_n_695);
  gl_ram_g13910 : AOI22D0BWP7T port map(A1 => gl_ram_ram_32(1), A2 => gl_ram_n_590, B1 => gl_ram_ram_35(1), B2 => gl_ram_n_584, ZN => gl_ram_n_694);
  gl_ram_g13911 : AOI22D0BWP7T port map(A1 => gl_ram_ram_9(2), A2 => gl_ram_n_588, B1 => gl_ram_ram_10(2), B2 => gl_ram_n_592, ZN => gl_ram_n_693);
  gl_ram_g13912 : AOI22D0BWP7T port map(A1 => gl_ram_ram_22(1), A2 => gl_ram_n_593, B1 => gl_ram_ram_23(1), B2 => gl_ram_n_587, ZN => gl_ram_n_692);
  gl_ram_g13913 : AOI22D0BWP7T port map(A1 => gl_ram_ram_84(1), A2 => gl_ram_n_586, B1 => gl_ram_ram_85(1), B2 => gl_ram_n_585, ZN => gl_ram_n_691);
  gl_ram_g13914 : AOI22D0BWP7T port map(A1 => gl_ram_ram_16(1), A2 => gl_ram_n_590, B1 => gl_ram_ram_19(1), B2 => gl_ram_n_584, ZN => gl_ram_n_690);
  gl_ram_g13915 : AOI22D0BWP7T port map(A1 => gl_ram_ram_12(2), A2 => gl_ram_n_586, B1 => gl_ram_ram_13(2), B2 => gl_ram_n_585, ZN => gl_ram_n_689);
  gl_ram_g13916 : AOI22D0BWP7T port map(A1 => gl_ram_ram_20(1), A2 => gl_ram_n_586, B1 => gl_ram_ram_21(1), B2 => gl_ram_n_585, ZN => gl_ram_n_688);
  gl_ram_g13917 : AOI22D0BWP7T port map(A1 => gl_ram_ram_49(2), A2 => gl_ram_n_588, B1 => gl_ram_ram_50(2), B2 => gl_ram_n_592, ZN => gl_ram_n_687);
  gl_ram_g13918 : AOI22D0BWP7T port map(A1 => FE_PHN511_gl_ram_ram_17_1, A2 => gl_ram_n_588, B1 => gl_ram_ram_18(1), B2 => gl_ram_n_592, ZN => gl_ram_n_686);
  gl_ram_g13919 : AOI22D0BWP7T port map(A1 => gl_ram_ram_70(2), A2 => gl_ram_n_593, B1 => gl_ram_ram_71(2), B2 => gl_ram_n_587, ZN => gl_ram_n_685);
  gl_ram_g13920 : AOI22D0BWP7T port map(A1 => gl_ram_ram_8(2), A2 => gl_ram_n_590, B1 => gl_ram_ram_11(2), B2 => gl_ram_n_584, ZN => gl_ram_n_684);
  gl_ram_g13921 : AOI22D0BWP7T port map(A1 => gl_ram_ram_25(0), A2 => gl_ram_n_588, B1 => gl_ram_ram_26(0), B2 => gl_ram_n_592, ZN => gl_ram_n_683);
  gl_ram_g13922 : AOI22D0BWP7T port map(A1 => gl_ram_ram_6(1), A2 => gl_ram_n_593, B1 => gl_ram_ram_7(1), B2 => gl_ram_n_587, ZN => gl_ram_n_682);
  gl_ram_g13923 : AOI22D0BWP7T port map(A1 => gl_ram_ram_1(1), A2 => gl_ram_n_588, B1 => gl_ram_ram_2(1), B2 => gl_ram_n_592, ZN => gl_ram_n_681);
  gl_ram_g13924 : AOI22D0BWP7T port map(A1 => gl_ram_ram_4(1), A2 => gl_ram_n_586, B1 => gl_ram_ram_5(1), B2 => gl_ram_n_585, ZN => gl_ram_n_680);
  gl_ram_g13925 : AOI22D0BWP7T port map(A1 => gl_ram_ram_22(2), A2 => gl_ram_n_593, B1 => gl_ram_ram_23(2), B2 => gl_ram_n_587, ZN => gl_ram_n_679);
  gl_ram_g13926 : AOI22D0BWP7T port map(A1 => gl_ram_ram_20(2), A2 => gl_ram_n_586, B1 => gl_ram_ram_21(2), B2 => gl_ram_n_585, ZN => gl_ram_n_678);
  gl_ram_g13927 : AOI22D0BWP7T port map(A1 => gl_ram_ram_0(1), A2 => gl_ram_n_590, B1 => gl_ram_ram_3(1), B2 => gl_ram_n_584, ZN => gl_ram_n_677);
  gl_ram_g13928 : AOI22D0BWP7T port map(A1 => gl_ram_ram_94(2), A2 => gl_ram_n_593, B1 => gl_ram_ram_95(2), B2 => gl_ram_n_587, ZN => gl_ram_n_676);
  gl_ram_g13929 : AOI22D0BWP7T port map(A1 => gl_ram_ram_65(2), A2 => gl_ram_n_588, B1 => gl_ram_ram_66(2), B2 => gl_ram_n_592, ZN => gl_ram_n_675);
  gl_ram_g13930 : AOI22D0BWP7T port map(A1 => gl_ram_ram_17(2), A2 => gl_ram_n_588, B1 => gl_ram_ram_18(2), B2 => gl_ram_n_592, ZN => gl_ram_n_674);
  gl_ram_g13931 : AOI22D0BWP7T port map(A1 => gl_ram_ram_68(2), A2 => gl_ram_n_586, B1 => gl_ram_ram_69(2), B2 => gl_ram_n_585, ZN => gl_ram_n_673);
  gl_ram_g13932 : AOI22D0BWP7T port map(A1 => gl_ram_ram_94(0), A2 => gl_ram_n_593, B1 => gl_ram_ram_95(0), B2 => gl_ram_n_587, ZN => gl_ram_n_672);
  gl_ram_g13933 : AOI22D0BWP7T port map(A1 => gl_ram_ram_16(2), A2 => gl_ram_n_590, B1 => gl_ram_ram_19(2), B2 => gl_ram_n_584, ZN => gl_ram_n_671);
  gl_ram_g13934 : AOI22D0BWP7T port map(A1 => gl_ram_ram_92(0), A2 => gl_ram_n_586, B1 => gl_ram_ram_93(0), B2 => gl_ram_n_585, ZN => gl_ram_n_670);
  gl_ram_g13935 : AOI22D0BWP7T port map(A1 => gl_ram_ram_89(0), A2 => gl_ram_n_588, B1 => gl_ram_ram_90(0), B2 => gl_ram_n_592, ZN => gl_ram_n_669);
  gl_ram_g13936 : AOI22D0BWP7T port map(A1 => gl_ram_ram_64(2), A2 => gl_ram_n_590, B1 => gl_ram_ram_67(2), B2 => gl_ram_n_584, ZN => gl_ram_n_668);
  gl_ram_g13937 : AOI22D0BWP7T port map(A1 => FE_PHN643_gl_ram_ram_88_0, A2 => gl_ram_n_590, B1 => gl_ram_ram_91(0), B2 => gl_ram_n_584, ZN => gl_ram_n_667);
  gl_ram_g13938 : AOI22D0BWP7T port map(A1 => gl_ram_ram_73(2), A2 => gl_ram_n_588, B1 => gl_ram_ram_74(2), B2 => gl_ram_n_592, ZN => gl_ram_n_666);
  gl_ram_g13939 : AOI22D0BWP7T port map(A1 => gl_ram_ram_64(1), A2 => gl_ram_n_590, B1 => gl_ram_ram_65(1), B2 => gl_ram_n_588, ZN => gl_ram_n_665);
  gl_ram_g13940 : AOI22D0BWP7T port map(A1 => gl_ram_ram_78(0), A2 => gl_ram_n_593, B1 => gl_ram_ram_79(0), B2 => gl_ram_n_587, ZN => gl_ram_n_664);
  gl_ram_g13941 : AOI22D0BWP7T port map(A1 => gl_ram_ram_72(0), A2 => gl_ram_n_590, B1 => gl_ram_ram_75(0), B2 => gl_ram_n_584, ZN => gl_ram_n_663);
  gl_ram_g13942 : AOI22D0BWP7T port map(A1 => gl_ram_ram_0(2), A2 => gl_ram_n_590, B1 => gl_ram_ram_3(2), B2 => gl_ram_n_584, ZN => gl_ram_n_662);
  gl_ram_g13943 : AOI22D0BWP7T port map(A1 => gl_ram_ram_76(0), A2 => gl_ram_n_586, B1 => gl_ram_ram_77(0), B2 => gl_ram_n_585, ZN => gl_ram_n_661);
  gl_ram_g13944 : AOI22D0BWP7T port map(A1 => gl_ram_ram_73(0), A2 => gl_ram_n_588, B1 => gl_ram_ram_74(0), B2 => gl_ram_n_592, ZN => gl_ram_n_660);
  gl_ram_g13945 : AOI22D0BWP7T port map(A1 => gl_ram_ram_4(2), A2 => gl_ram_n_586, B1 => gl_ram_ram_5(2), B2 => gl_ram_n_585, ZN => gl_ram_n_659);
  gl_ram_g13946 : AOI22D0BWP7T port map(A1 => gl_ram_ram_86(0), A2 => gl_ram_n_593, B1 => gl_ram_ram_87(0), B2 => gl_ram_n_587, ZN => gl_ram_n_658);
  gl_ram_g13947 : AOI22D0BWP7T port map(A1 => gl_ram_ram_1(2), A2 => gl_ram_n_588, B1 => gl_ram_ram_2(2), B2 => gl_ram_n_592, ZN => gl_ram_n_657);
  gl_ram_g13948 : AOI22D0BWP7T port map(A1 => gl_ram_ram_81(0), A2 => gl_ram_n_588, B1 => gl_ram_ram_82(0), B2 => gl_ram_n_592, ZN => gl_ram_n_656);
  gl_ram_g13949 : AOI22D0BWP7T port map(A1 => gl_ram_ram_84(0), A2 => gl_ram_n_586, B1 => gl_ram_ram_85(0), B2 => gl_ram_n_585, ZN => gl_ram_n_655);
  gl_ram_g13950 : AOI22D0BWP7T port map(A1 => gl_ram_ram_80(0), A2 => gl_ram_n_590, B1 => gl_ram_ram_83(0), B2 => gl_ram_n_584, ZN => gl_ram_n_654);
  gl_ram_g13951 : AOI22D0BWP7T port map(A1 => gl_ram_ram_62(2), A2 => gl_ram_n_593, B1 => gl_ram_ram_63(2), B2 => gl_ram_n_587, ZN => gl_ram_n_653);
  gl_ram_g13952 : AOI22D0BWP7T port map(A1 => gl_ram_ram_70(0), A2 => gl_ram_n_593, B1 => gl_ram_ram_71(0), B2 => gl_ram_n_587, ZN => gl_ram_n_652);
  gl_ram_g13953 : AOI22D0BWP7T port map(A1 => gl_ram_ram_92(2), A2 => gl_ram_n_586, B1 => gl_ram_ram_93(2), B2 => gl_ram_n_585, ZN => gl_ram_n_651);
  gl_ram_g13954 : AOI22D0BWP7T port map(A1 => gl_ram_ram_64(0), A2 => gl_ram_n_590, B1 => gl_ram_ram_67(0), B2 => gl_ram_n_584, ZN => gl_ram_n_650);
  gl_ram_g13955 : AOI22D0BWP7T port map(A1 => gl_ram_ram_68(0), A2 => gl_ram_n_586, B1 => gl_ram_ram_69(0), B2 => gl_ram_n_585, ZN => gl_ram_n_649);
  gl_ram_g13956 : AOI22D0BWP7T port map(A1 => gl_ram_ram_65(0), A2 => gl_ram_n_588, B1 => gl_ram_ram_66(0), B2 => gl_ram_n_592, ZN => gl_ram_n_648);
  gl_ram_g13957 : AOI22D0BWP7T port map(A1 => gl_ram_ram_57(2), A2 => gl_ram_n_588, B1 => gl_ram_ram_58(2), B2 => gl_ram_n_592, ZN => gl_ram_n_647);
  gl_ram_g13958 : AOI22D0BWP7T port map(A1 => gl_ram_ram_62(0), A2 => gl_ram_n_593, B1 => gl_ram_ram_63(0), B2 => gl_ram_n_587, ZN => gl_ram_n_646);
  gl_ram_g13959 : AOI22D0BWP7T port map(A1 => gl_ram_ram_94(1), A2 => gl_ram_n_593, B1 => gl_ram_ram_95(1), B2 => gl_ram_n_587, ZN => gl_ram_n_645);
  gl_ram_g13960 : AOI22D0BWP7T port map(A1 => gl_ram_ram_60(0), A2 => gl_ram_n_586, B1 => gl_ram_ram_61(0), B2 => gl_ram_n_585, ZN => gl_ram_n_644);
  gl_ram_g13961 : AOI22D0BWP7T port map(A1 => gl_ram_ram_60(2), A2 => gl_ram_n_586, B1 => gl_ram_ram_61(2), B2 => gl_ram_n_585, ZN => gl_ram_n_643);
  gl_ram_g13962 : AOI22D0BWP7T port map(A1 => gl_ram_ram_89(1), A2 => gl_ram_n_588, B1 => gl_ram_ram_90(1), B2 => gl_ram_n_592, ZN => gl_ram_n_642);
  gl_ram_g13963 : AOI22D0BWP7T port map(A1 => gl_ram_ram_57(0), A2 => gl_ram_n_588, B1 => gl_ram_ram_58(0), B2 => gl_ram_n_592, ZN => gl_ram_n_641);
  gl_ram_g13964 : AOI22D0BWP7T port map(A1 => gl_ram_ram_56(0), A2 => gl_ram_n_590, B1 => gl_ram_ram_59(0), B2 => gl_ram_n_584, ZN => gl_ram_n_640);
  gl_ram_g13965 : AOI22D0BWP7T port map(A1 => gl_ram_ram_92(1), A2 => gl_ram_n_586, B1 => gl_ram_ram_93(1), B2 => gl_ram_n_585, ZN => gl_ram_n_639);
  gl_ram_g13966 : AOI22D0BWP7T port map(A1 => gl_ram_ram_54(0), A2 => gl_ram_n_593, B1 => gl_ram_ram_55(0), B2 => gl_ram_n_587, ZN => gl_ram_n_638);
  gl_ram_g13967 : AOI22D0BWP7T port map(A1 => gl_ram_ram_49(0), A2 => gl_ram_n_588, B1 => gl_ram_ram_50(0), B2 => gl_ram_n_592, ZN => gl_ram_n_637);
  gl_ram_g13968 : AOI22D0BWP7T port map(A1 => gl_ram_ram_88(1), A2 => gl_ram_n_590, B1 => gl_ram_ram_91(1), B2 => gl_ram_n_584, ZN => gl_ram_n_636);
  gl_ram_g13969 : AOI22D0BWP7T port map(A1 => gl_ram_ram_56(2), A2 => gl_ram_n_590, B1 => gl_ram_ram_59(2), B2 => gl_ram_n_584, ZN => gl_ram_n_635);
  gl_ram_g13970 : AOI22D0BWP7T port map(A1 => gl_ram_ram_52(0), A2 => gl_ram_n_586, B1 => gl_ram_ram_53(0), B2 => gl_ram_n_585, ZN => gl_ram_n_634);
  gl_ram_g13971 : AOI22D0BWP7T port map(A1 => gl_ram_ram_48(0), A2 => gl_ram_n_590, B1 => gl_ram_ram_51(0), B2 => gl_ram_n_584, ZN => gl_ram_n_633);
  gl_ram_g13972 : AOI22D0BWP7T port map(A1 => gl_ram_ram_89(2), A2 => gl_ram_n_588, B1 => gl_ram_ram_90(2), B2 => gl_ram_n_592, ZN => gl_ram_n_632);
  gl_ram_g13973 : AOI22D0BWP7T port map(A1 => gl_ram_ram_46(0), A2 => gl_ram_n_593, B1 => gl_ram_ram_47(0), B2 => gl_ram_n_587, ZN => gl_ram_n_631);
  gl_ram_g13974 : AOI22D0BWP7T port map(A1 => gl_ram_ram_78(1), A2 => gl_ram_n_593, B1 => gl_ram_ram_79(1), B2 => gl_ram_n_587, ZN => gl_ram_n_630);
  gl_ram_g13975 : AOI22D0BWP7T port map(A1 => gl_ram_ram_41(0), A2 => gl_ram_n_588, B1 => gl_ram_ram_42(0), B2 => gl_ram_n_592, ZN => gl_ram_n_629);
  gl_ram_g13976 : AOI22D0BWP7T port map(A1 => gl_ram_ram_72(1), A2 => gl_ram_n_590, B1 => gl_ram_ram_75(1), B2 => gl_ram_n_584, ZN => gl_ram_n_628);
  gl_ram_g13977 : AOI22D0BWP7T port map(A1 => gl_ram_ram_44(0), A2 => gl_ram_n_586, B1 => gl_ram_ram_45(0), B2 => gl_ram_n_585, ZN => gl_ram_n_627);
  gl_ram_g13978 : AOI22D0BWP7T port map(A1 => gl_ram_ram_40(0), A2 => gl_ram_n_590, B1 => gl_ram_ram_43(0), B2 => gl_ram_n_584, ZN => gl_ram_n_626);
  gl_ram_g13979 : AOI22D0BWP7T port map(A1 => gl_ram_ram_54(2), A2 => gl_ram_n_593, B1 => gl_ram_ram_55(2), B2 => gl_ram_n_587, ZN => gl_ram_n_625);
  gl_ram_g13980 : AOI22D0BWP7T port map(A1 => gl_ram_ram_76(1), A2 => gl_ram_n_586, B1 => gl_ram_ram_77(1), B2 => gl_ram_n_585, ZN => gl_ram_n_624);
  gl_ram_g13981 : AOI22D0BWP7T port map(A1 => gl_ram_ram_38(0), A2 => gl_ram_n_593, B1 => gl_ram_ram_39(0), B2 => gl_ram_n_587, ZN => gl_ram_n_623);
  gl_ram_g13982 : AOI22D0BWP7T port map(A1 => gl_ram_ram_73(1), A2 => gl_ram_n_588, B1 => gl_ram_ram_74(1), B2 => gl_ram_n_592, ZN => gl_ram_n_622);
  gl_ram_g13983 : AOI22D0BWP7T port map(A1 => gl_ram_ram_33(0), A2 => gl_ram_n_588, B1 => gl_ram_ram_34(0), B2 => gl_ram_n_592, ZN => gl_ram_n_621);
  gl_ram_g13984 : AOI22D0BWP7T port map(A1 => gl_ram_ram_36(0), A2 => gl_ram_n_586, B1 => gl_ram_ram_37(0), B2 => gl_ram_n_585, ZN => gl_ram_n_620);
  gl_ram_g13985 : AOI22D0BWP7T port map(A1 => gl_ram_ram_32(0), A2 => gl_ram_n_590, B1 => gl_ram_ram_35(0), B2 => gl_ram_n_584, ZN => gl_ram_n_619);
  gl_ram_g13986 : AOI22D0BWP7T port map(A1 => gl_ram_ram_48(2), A2 => gl_ram_n_590, B1 => gl_ram_ram_51(2), B2 => gl_ram_n_584, ZN => gl_ram_n_618);
  gl_ram_g13987 : AOI22D0BWP7T port map(A1 => gl_ram_ram_86(1), A2 => gl_ram_n_593, B1 => gl_ram_ram_87(1), B2 => gl_ram_n_587, ZN => gl_ram_n_617);
  gl_ram_g13988 : AOI22D0BWP7T port map(A1 => gl_ram_ram_30(0), A2 => gl_ram_n_593, B1 => gl_ram_ram_31(0), B2 => gl_ram_n_587, ZN => gl_ram_n_616);
  gl_ram_g13989 : AOI22D0BWP7T port map(A1 => gl_ram_ram_28(0), A2 => gl_ram_n_586, B1 => gl_ram_ram_29(0), B2 => gl_ram_n_585, ZN => gl_ram_n_615);
  gl_ram_g13990 : AOI22D0BWP7T port map(A1 => gl_ram_ram_81(1), A2 => gl_ram_n_588, B1 => gl_ram_ram_82(1), B2 => gl_ram_n_592, ZN => gl_ram_n_614);
  gl_ram_g13991 : AOI22D0BWP7T port map(A1 => gl_ram_ram_24(0), A2 => gl_ram_n_590, B1 => gl_ram_ram_27(0), B2 => gl_ram_n_584, ZN => gl_ram_n_613);
  gl_ram_g13992 : AOI22D0BWP7T port map(A1 => gl_ram_ram_52(2), A2 => gl_ram_n_586, B1 => gl_ram_ram_53(2), B2 => gl_ram_n_585, ZN => gl_ram_n_612);
  gl_ram_g13993 : AOI22D0BWP7T port map(A1 => gl_ram_ram_14(0), A2 => gl_ram_n_593, B1 => gl_ram_ram_15(0), B2 => gl_ram_n_587, ZN => gl_ram_n_611);
  gl_ram_g13994 : AOI22D0BWP7T port map(A1 => gl_ram_ram_8(0), A2 => gl_ram_n_590, B1 => gl_ram_ram_11(0), B2 => gl_ram_n_584, ZN => gl_ram_n_610);
  gl_ram_g13995 : AOI22D0BWP7T port map(A1 => gl_ram_ram_80(1), A2 => gl_ram_n_590, B1 => gl_ram_ram_83(1), B2 => gl_ram_n_584, ZN => gl_ram_n_609);
  gl_ram_g13996 : AOI22D0BWP7T port map(A1 => gl_ram_ram_12(0), A2 => gl_ram_n_586, B1 => gl_ram_ram_13(0), B2 => gl_ram_n_585, ZN => gl_ram_n_608);
  gl_ram_g13997 : AOI22D0BWP7T port map(A1 => gl_ram_ram_9(0), A2 => gl_ram_n_588, B1 => gl_ram_ram_10(0), B2 => gl_ram_n_592, ZN => gl_ram_n_607);
  gl_ram_g13998 : AOI22D0BWP7T port map(A1 => gl_ram_ram_70(1), A2 => gl_ram_n_593, B1 => gl_ram_ram_71(1), B2 => gl_ram_n_587, ZN => gl_ram_n_606);
  gl_ram_g13999 : AOI22D0BWP7T port map(A1 => gl_ram_ram_22(0), A2 => gl_ram_n_593, B1 => gl_ram_ram_23(0), B2 => gl_ram_n_587, ZN => gl_ram_n_605);
  gl_ram_g14000 : AOI22D0BWP7T port map(A1 => gl_ram_ram_20(0), A2 => gl_ram_n_586, B1 => gl_ram_ram_21(0), B2 => gl_ram_n_585, ZN => gl_ram_n_604);
  gl_ram_g14001 : AOI22D0BWP7T port map(A1 => gl_ram_ram_76(2), A2 => gl_ram_n_586, B1 => gl_ram_ram_77(2), B2 => gl_ram_n_585, ZN => gl_ram_n_603);
  gl_ram_g14002 : AOI22D0BWP7T port map(A1 => gl_ram_ram_68(1), A2 => gl_ram_n_586, B1 => gl_ram_ram_69(1), B2 => gl_ram_n_585, ZN => gl_ram_n_602);
  gl_ram_g14003 : AOI22D0BWP7T port map(A1 => gl_ram_ram_18(0), A2 => gl_ram_n_592, B1 => gl_ram_ram_19(0), B2 => gl_ram_n_584, ZN => gl_ram_n_601);
  gl_ram_g14004 : AOI22D0BWP7T port map(A1 => gl_ram_ram_16(0), A2 => gl_ram_n_590, B1 => gl_ram_ram_17(0), B2 => gl_ram_n_588, ZN => gl_ram_n_600);
  gl_ram_g14005 : AOI22D0BWP7T port map(A1 => gl_ram_ram_6(0), A2 => gl_ram_n_593, B1 => gl_ram_ram_7(0), B2 => gl_ram_n_587, ZN => gl_ram_n_599);
  gl_ram_g14006 : AOI22D0BWP7T port map(A1 => gl_ram_ram_46(2), A2 => gl_ram_n_593, B1 => gl_ram_ram_47(2), B2 => gl_ram_n_587, ZN => gl_ram_n_598);
  gl_ram_g14007 : AOI22D0BWP7T port map(A1 => gl_ram_ram_0(0), A2 => gl_ram_n_590, B1 => gl_ram_ram_3(0), B2 => gl_ram_n_584, ZN => gl_ram_n_597);
  gl_ram_g14008 : AOI22D0BWP7T port map(A1 => gl_ram_ram_4(0), A2 => gl_ram_n_586, B1 => gl_ram_ram_5(0), B2 => gl_ram_n_585, ZN => gl_ram_n_596);
  gl_ram_g14009 : AOI22D0BWP7T port map(A1 => gl_ram_ram_1(0), A2 => gl_ram_n_588, B1 => gl_ram_ram_2(0), B2 => gl_ram_n_592, ZN => gl_ram_n_595);
  gl_ram_g14010 : AOI22D0BWP7T port map(A1 => gl_ram_ram_6(2), A2 => gl_ram_n_593, B1 => gl_ram_ram_7(2), B2 => gl_ram_n_587, ZN => gl_ram_n_594);
  gl_ram_g14011 : INVD1BWP7T port map(I => gl_ram_n_591, ZN => gl_ram_n_592);
  gl_ram_g14012 : INVD1BWP7T port map(I => gl_ram_n_589, ZN => gl_ram_n_590);
  gl_ram_g14014 : AN2D1BWP7T port map(A1 => gl_ram_n_583, A2 => gl_ram_n_579, Z => gl_ram_n_593);
  gl_ram_g14015 : ND2D0BWP7T port map(A1 => gl_ram_n_582, A2 => gl_ram_n_579, ZN => gl_ram_n_591);
  gl_ram_g14016 : ND2D0BWP7T port map(A1 => gl_ram_n_582, A2 => gl_ram_n_577, ZN => gl_ram_n_589);
  gl_ram_g14017 : NR2XD1BWP7T port map(A1 => gl_ram_n_583, A2 => gl_ram_n_580, ZN => gl_ram_n_588);
  gl_ram_g14019 : NR2XD1BWP7T port map(A1 => gl_ram_n_582, A2 => gl_ram_n_578, ZN => gl_ram_n_587);
  gl_ram_g14020 : AN2D1BWP7T port map(A1 => gl_ram_n_583, A2 => gl_ram_n_577, Z => gl_ram_n_586);
  gl_ram_g14021 : NR2XD1BWP7T port map(A1 => gl_ram_n_582, A2 => gl_ram_n_580, ZN => gl_ram_n_585);
  gl_ram_g14022 : NR2XD1BWP7T port map(A1 => gl_ram_n_583, A2 => gl_ram_n_578, ZN => gl_ram_n_584);
  gl_ram_g14023 : INVD1BWP7T port map(I => gl_ram_n_583, ZN => gl_ram_n_582);
  gl_ram_g14024 : FA1D0BWP7T port map(A => gl_sig_x(2), B => gl_sig_y(1), CI => gl_ram_n_571, CO => gl_ram_n_581, S => gl_ram_n_583);
  gl_ram_g14025 : ND2D0BWP7T port map(A1 => gl_ram_n_572, A2 => gl_sig_x(0), ZN => gl_ram_n_580);
  gl_ram_g14026 : NR2D0BWP7T port map(A1 => gl_ram_n_572, A2 => gl_sig_x(0), ZN => gl_ram_n_579);
  gl_ram_g14027 : IND2D0BWP7T port map(A1 => gl_ram_n_572, B1 => gl_sig_x(0), ZN => gl_ram_n_578);
  gl_ram_g14028 : INR2D0BWP7T port map(A1 => gl_ram_n_572, B1 => gl_sig_x(0), ZN => gl_ram_n_577);
  gl_ram_g14029 : HA1D0BWP7T port map(A => gl_sig_x(3), B => gl_sig_y(0), CO => gl_ram_n_575, S => gl_ram_n_576);
  gl_ram_g14030 : HA1D0BWP7T port map(A => gl_sig_y(3), B => gl_sig_y(1), CO => gl_ram_n_573, S => gl_ram_n_574);
  gl_ram_g14031 : XNR2D1BWP7T port map(A1 => gl_sig_y(0), A2 => gl_sig_x(1), ZN => gl_ram_n_572);
  gl_ram_g14032 : AN2D1BWP7T port map(A1 => gl_sig_y(0), A2 => gl_sig_x(1), Z => gl_ram_n_571);
  gl_ram_g2 : INR2D1BWP7T port map(A1 => gl_ram_n_588, B1 => gl_ram_n_790, ZN => gl_ram_n_570);
  gl_ram_g14033 : INR2D1BWP7T port map(A1 => gl_ram_n_584, B1 => gl_ram_n_790, ZN => gl_ram_n_569);
  gl_ram_ram_position_reg_0 : DFQD1BWP7T port map(CP => CTS_19, D => FE_PHN360_gl_ram_n_142, Q => gl_ram_ram_position(0));
  gl_ram_ram_position_reg_1 : DFQD1BWP7T port map(CP => CTS_19, D => FE_PHN376_gl_ram_n_308, Q => gl_ram_ram_position(1));
  gl_ram_ram_position_reg_2 : DFQD1BWP7T port map(CP => CTS_23, D => FE_PHN375_gl_ram_n_552, Q => gl_ram_ram_position(2));
  gl_ram_ram_position_reg_3 : DFQD1BWP7T port map(CP => CTS_23, D => FE_PHN389_gl_ram_n_563, Q => gl_ram_ram_position(3));
  gl_ram_ram_position_reg_5 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_567, Q => gl_ram_ram_position(5));
  gl_ram_ram_position_reg_6 : DFQD1BWP7T port map(CP => CTS_23, D => FE_PHN382_gl_ram_n_564, Q => gl_ram_ram_position(6));
  gl_ram_ram_reg_0_0 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_356, Q => gl_ram_ram_0(0));
  gl_ram_ram_reg_0_1 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_351, Q => gl_ram_ram_0(1));
  gl_ram_ram_reg_0_2 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_330, Q => gl_ram_ram_0(2));
  gl_ram_ram_reg_1_0 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_321, Q => gl_ram_ram_1(0));
  gl_ram_ram_reg_1_1 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_533, Q => gl_ram_ram_1(1));
  gl_ram_ram_reg_1_2 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_551, Q => gl_ram_ram_1(2));
  gl_ram_ram_reg_2_0 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_538, Q => gl_ram_ram_2(0));
  gl_ram_ram_reg_2_1 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_532, Q => gl_ram_ram_2(1));
  gl_ram_ram_reg_2_2 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_529, Q => gl_ram_ram_2(2));
  gl_ram_ram_reg_3_0 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_526, Q => gl_ram_ram_3(0));
  gl_ram_ram_reg_3_1 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_519, Q => gl_ram_ram_3(1));
  gl_ram_ram_reg_3_2 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_517, Q => gl_ram_ram_3(2));
  gl_ram_ram_reg_4_0 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_514, Q => gl_ram_ram_4(0));
  gl_ram_ram_reg_4_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_509, Q => gl_ram_ram_4(1));
  gl_ram_ram_reg_4_2 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_508, Q => gl_ram_ram_4(2));
  gl_ram_ram_reg_5_0 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_503, Q => gl_ram_ram_5(0));
  gl_ram_ram_reg_5_1 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_498, Q => gl_ram_ram_5(1));
  gl_ram_ram_reg_5_2 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_491, Q => gl_ram_ram_5(2));
  gl_ram_ram_reg_6_0 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_493, Q => gl_ram_ram_6(0));
  gl_ram_ram_reg_6_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_486, Q => gl_ram_ram_6(1));
  gl_ram_ram_reg_6_2 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_485, Q => gl_ram_ram_6(2));
  gl_ram_ram_reg_7_0 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_481, Q => gl_ram_ram_7(0));
  gl_ram_ram_reg_7_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_479, Q => gl_ram_ram_7(1));
  gl_ram_ram_reg_7_2 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_474, Q => gl_ram_ram_7(2));
  gl_ram_ram_reg_8_0 : DFQD1BWP7T port map(CP => CTS_22, D => FE_PHN672_gl_ram_n_470, Q => gl_ram_ram_8(0));
  gl_ram_ram_reg_8_1 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_467, Q => FE_PHN647_gl_ram_ram_8_1);
  gl_ram_ram_reg_8_2 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_554, Q => gl_ram_ram_8(2));
  gl_ram_ram_reg_9_0 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_458, Q => gl_ram_ram_9(0));
  gl_ram_ram_reg_9_1 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_461, Q => gl_ram_ram_9(1));
  gl_ram_ram_reg_9_2 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_457, Q => gl_ram_ram_9(2));
  gl_ram_ram_reg_10_0 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_454, Q => gl_ram_ram_10(0));
  gl_ram_ram_reg_10_1 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_451, Q => gl_ram_ram_10(1));
  gl_ram_ram_reg_10_2 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_448, Q => gl_ram_ram_10(2));
  gl_ram_ram_reg_11_0 : DFQD1BWP7T port map(CP => CTS_22, D => FE_PHN657_gl_ram_n_445, Q => gl_ram_ram_11(0));
  gl_ram_ram_reg_11_1 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_442, Q => gl_ram_ram_11(1));
  gl_ram_ram_reg_11_2 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_439, Q => FE_PHN652_gl_ram_ram_11_2);
  gl_ram_ram_reg_12_0 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_436, Q => gl_ram_ram_12(0));
  gl_ram_ram_reg_12_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_433, Q => FE_PHN642_gl_ram_ram_12_1);
  gl_ram_ram_reg_12_2 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_430, Q => gl_ram_ram_12(2));
  gl_ram_ram_reg_13_0 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_428, Q => gl_ram_ram_13(0));
  gl_ram_ram_reg_13_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_424, Q => gl_ram_ram_13(1));
  gl_ram_ram_reg_13_2 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_421, Q => gl_ram_ram_13(2));
  gl_ram_ram_reg_14_0 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_418, Q => gl_ram_ram_14(0));
  gl_ram_ram_reg_14_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_415, Q => gl_ram_ram_14(1));
  gl_ram_ram_reg_14_2 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_412, Q => gl_ram_ram_14(2));
  gl_ram_ram_reg_15_0 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_410, Q => gl_ram_ram_15(0));
  gl_ram_ram_reg_15_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_406, Q => gl_ram_ram_15(1));
  gl_ram_ram_reg_15_2 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_403, Q => gl_ram_ram_15(2));
  gl_ram_ram_reg_16_0 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_402, Q => gl_ram_ram_16(0));
  gl_ram_ram_reg_16_1 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_401, Q => gl_ram_ram_16(1));
  gl_ram_ram_reg_16_2 : DFQD1BWP7T port map(CP => CTS_22, D => FE_PHN469_gl_ram_n_400, Q => FE_PHN651_gl_ram_ram_16_2);
  gl_ram_ram_reg_17_0 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_399, Q => gl_ram_ram_17(0));
  gl_ram_ram_reg_17_1 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_398, Q => gl_ram_ram_17(1));
  gl_ram_ram_reg_17_2 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_397, Q => gl_ram_ram_17(2));
  gl_ram_ram_reg_18_0 : DFQD1BWP7T port map(CP => CTS_22, D => FE_PHN471_gl_ram_n_396, Q => gl_ram_ram_18(0));
  gl_ram_ram_reg_18_1 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_395, Q => gl_ram_ram_18(1));
  gl_ram_ram_reg_18_2 : DFQD1BWP7T port map(CP => CTS_22, D => FE_PHN413_gl_ram_n_394, Q => gl_ram_ram_18(2));
  gl_ram_ram_reg_19_0 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_393, Q => gl_ram_ram_19(0));
  gl_ram_ram_reg_19_1 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_392, Q => FE_PHN611_gl_ram_ram_19_1);
  gl_ram_ram_reg_19_2 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_391, Q => gl_ram_ram_19(2));
  gl_ram_ram_reg_20_0 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_390, Q => gl_ram_ram_20(0));
  gl_ram_ram_reg_20_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_389, Q => gl_ram_ram_20(1));
  gl_ram_ram_reg_20_2 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_388, Q => gl_ram_ram_20(2));
  gl_ram_ram_reg_21_0 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_387, Q => gl_ram_ram_21(0));
  gl_ram_ram_reg_21_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_386, Q => gl_ram_ram_21(1));
  gl_ram_ram_reg_21_2 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_385, Q => gl_ram_ram_21(2));
  gl_ram_ram_reg_22_0 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_384, Q => gl_ram_ram_22(0));
  gl_ram_ram_reg_22_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_383, Q => gl_ram_ram_22(1));
  gl_ram_ram_reg_22_2 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_382, Q => gl_ram_ram_22(2));
  gl_ram_ram_reg_23_0 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_381, Q => gl_ram_ram_23(0));
  gl_ram_ram_reg_23_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_380, Q => gl_ram_ram_23(1));
  gl_ram_ram_reg_23_2 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_379, Q => gl_ram_ram_23(2));
  gl_ram_ram_reg_24_0 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_377, Q => gl_ram_ram_24(0));
  gl_ram_ram_reg_24_1 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_373, Q => gl_ram_ram_24(1));
  gl_ram_ram_reg_24_2 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_370, Q => gl_ram_ram_24(2));
  gl_ram_ram_reg_25_0 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_367, Q => gl_ram_ram_25(0));
  gl_ram_ram_reg_25_1 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_364, Q => gl_ram_ram_25(1));
  gl_ram_ram_reg_25_2 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_361, Q => gl_ram_ram_25(2));
  gl_ram_ram_reg_26_0 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_358, Q => gl_ram_ram_26(0));
  gl_ram_ram_reg_26_1 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_354, Q => gl_ram_ram_26(1));
  gl_ram_ram_reg_26_2 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_349, Q => gl_ram_ram_26(2));
  gl_ram_ram_reg_27_0 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_347, Q => gl_ram_ram_27(0));
  gl_ram_ram_reg_27_1 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_344, Q => gl_ram_ram_27(1));
  gl_ram_ram_reg_27_2 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_340, Q => FE_PHN669_gl_ram_ram_27_2);
  gl_ram_ram_reg_28_0 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_338, Q => gl_ram_ram_28(0));
  gl_ram_ram_reg_28_1 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_335, Q => gl_ram_ram_28(1));
  gl_ram_ram_reg_28_2 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_332, Q => gl_ram_ram_28(2));
  gl_ram_ram_reg_29_0 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_328, Q => gl_ram_ram_29(0));
  gl_ram_ram_reg_29_1 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_325, Q => gl_ram_ram_29(1));
  gl_ram_ram_reg_29_2 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_323, Q => gl_ram_ram_29(2));
  gl_ram_ram_reg_30_0 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_318, Q => gl_ram_ram_30(0));
  gl_ram_ram_reg_30_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_315, Q => gl_ram_ram_30(1));
  gl_ram_ram_reg_30_2 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_548, Q => gl_ram_ram_30(2));
  gl_ram_ram_reg_31_0 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_546, Q => gl_ram_ram_31(0));
  gl_ram_ram_reg_31_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_543, Q => gl_ram_ram_31(1));
  gl_ram_ram_reg_31_2 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_540, Q => gl_ram_ram_31(2));
  gl_ram_ram_reg_32_0 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_539, Q => gl_ram_ram_32(0));
  gl_ram_ram_reg_32_1 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_536, Q => gl_ram_ram_32(1));
  gl_ram_ram_reg_32_2 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_537, Q => gl_ram_ram_32(2));
  gl_ram_ram_reg_33_0 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_535, Q => gl_ram_ram_33(0));
  gl_ram_ram_reg_33_1 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_534, Q => gl_ram_ram_33(1));
  gl_ram_ram_reg_33_2 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_531, Q => gl_ram_ram_33(2));
  gl_ram_ram_reg_34_0 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_530, Q => gl_ram_ram_34(0));
  gl_ram_ram_reg_34_1 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_528, Q => gl_ram_ram_34(1));
  gl_ram_ram_reg_34_2 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_527, Q => gl_ram_ram_34(2));
  gl_ram_ram_reg_35_0 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_525, Q => gl_ram_ram_35(0));
  gl_ram_ram_reg_35_1 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_524, Q => gl_ram_ram_35(1));
  gl_ram_ram_reg_35_2 : DFQD1BWP7T port map(CP => CTS_22, D => FE_PHN627_gl_ram_n_523, Q => gl_ram_ram_35(2));
  gl_ram_ram_reg_36_0 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_522, Q => gl_ram_ram_36(0));
  gl_ram_ram_reg_36_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_521, Q => gl_ram_ram_36(1));
  gl_ram_ram_reg_36_2 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_520, Q => gl_ram_ram_36(2));
  gl_ram_ram_reg_37_0 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_518, Q => gl_ram_ram_37(0));
  gl_ram_ram_reg_37_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_516, Q => gl_ram_ram_37(1));
  gl_ram_ram_reg_37_2 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_515, Q => gl_ram_ram_37(2));
  gl_ram_ram_reg_38_0 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_513, Q => gl_ram_ram_38(0));
  gl_ram_ram_reg_38_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_512, Q => gl_ram_ram_38(1));
  gl_ram_ram_reg_38_2 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_511, Q => gl_ram_ram_38(2));
  gl_ram_ram_reg_39_0 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_510, Q => gl_ram_ram_39(0));
  gl_ram_ram_reg_39_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_507, Q => gl_ram_ram_39(1));
  gl_ram_ram_reg_39_2 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_506, Q => gl_ram_ram_39(2));
  gl_ram_ram_reg_40_0 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_505, Q => gl_ram_ram_40(0));
  gl_ram_ram_reg_40_1 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_504, Q => gl_ram_ram_40(1));
  gl_ram_ram_reg_40_2 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_502, Q => gl_ram_ram_40(2));
  gl_ram_ram_reg_41_0 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_501, Q => gl_ram_ram_41(0));
  gl_ram_ram_reg_41_1 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_500, Q => gl_ram_ram_41(1));
  gl_ram_ram_reg_41_2 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_499, Q => gl_ram_ram_41(2));
  gl_ram_ram_reg_42_0 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_497, Q => gl_ram_ram_42(0));
  gl_ram_ram_reg_42_1 : DFQD1BWP7T port map(CP => CTS_22, D => FE_PHN415_gl_ram_n_496, Q => gl_ram_ram_42(1));
  gl_ram_ram_reg_42_2 : DFQD1BWP7T port map(CP => CTS_22, D => FE_PHN425_gl_ram_n_495, Q => gl_ram_ram_42(2));
  gl_ram_ram_reg_43_0 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_494, Q => gl_ram_ram_43(0));
  gl_ram_ram_reg_43_1 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_492, Q => gl_ram_ram_43(1));
  gl_ram_ram_reg_43_2 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_490, Q => gl_ram_ram_43(2));
  gl_ram_ram_reg_44_0 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_489, Q => gl_ram_ram_44(0));
  gl_ram_ram_reg_44_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_488, Q => gl_ram_ram_44(1));
  gl_ram_ram_reg_44_2 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_487, Q => gl_ram_ram_44(2));
  gl_ram_ram_reg_45_0 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_484, Q => gl_ram_ram_45(0));
  gl_ram_ram_reg_45_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_483, Q => gl_ram_ram_45(1));
  gl_ram_ram_reg_45_2 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_482, Q => gl_ram_ram_45(2));
  gl_ram_ram_reg_46_0 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_480, Q => gl_ram_ram_46(0));
  gl_ram_ram_reg_46_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_478, Q => gl_ram_ram_46(1));
  gl_ram_ram_reg_46_2 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_477, Q => gl_ram_ram_46(2));
  gl_ram_ram_reg_47_0 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_476, Q => gl_ram_ram_47(0));
  gl_ram_ram_reg_47_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_475, Q => gl_ram_ram_47(1));
  gl_ram_ram_reg_47_2 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_473, Q => gl_ram_ram_47(2));
  gl_ram_ram_reg_48_0 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_472, Q => gl_ram_ram_48(0));
  gl_ram_ram_reg_48_1 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_471, Q => gl_ram_ram_48(1));
  gl_ram_ram_reg_48_2 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_469, Q => gl_ram_ram_48(2));
  gl_ram_ram_reg_49_0 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_468, Q => gl_ram_ram_49(0));
  gl_ram_ram_reg_49_1 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_466, Q => gl_ram_ram_49(1));
  gl_ram_ram_reg_49_2 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_465, Q => gl_ram_ram_49(2));
  gl_ram_ram_reg_50_0 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_553, Q => gl_ram_ram_50(0));
  gl_ram_ram_reg_50_1 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_464, Q => gl_ram_ram_50(1));
  gl_ram_ram_reg_50_2 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_463, Q => gl_ram_ram_50(2));
  gl_ram_ram_reg_51_0 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_462, Q => gl_ram_ram_51(0));
  gl_ram_ram_reg_51_1 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_460, Q => gl_ram_ram_51(1));
  gl_ram_ram_reg_51_2 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_459, Q => gl_ram_ram_51(2));
  gl_ram_ram_reg_52_0 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_456, Q => gl_ram_ram_52(0));
  gl_ram_ram_reg_52_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_455, Q => gl_ram_ram_52(1));
  gl_ram_ram_reg_52_2 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_453, Q => gl_ram_ram_52(2));
  gl_ram_ram_reg_53_0 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_452, Q => gl_ram_ram_53(0));
  gl_ram_ram_reg_53_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_450, Q => gl_ram_ram_53(1));
  gl_ram_ram_reg_53_2 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_449, Q => gl_ram_ram_53(2));
  gl_ram_ram_reg_54_0 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_447, Q => gl_ram_ram_54(0));
  gl_ram_ram_reg_54_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_446, Q => gl_ram_ram_54(1));
  gl_ram_ram_reg_54_2 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_444, Q => gl_ram_ram_54(2));
  gl_ram_ram_reg_55_0 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_443, Q => gl_ram_ram_55(0));
  gl_ram_ram_reg_55_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_441, Q => gl_ram_ram_55(1));
  gl_ram_ram_reg_55_2 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_440, Q => gl_ram_ram_55(2));
  gl_ram_ram_reg_56_0 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_438, Q => gl_ram_ram_56(0));
  gl_ram_ram_reg_56_1 : DFQD1BWP7T port map(CP => CTS_21, D => FE_PHN628_gl_ram_n_437, Q => gl_ram_ram_56(1));
  gl_ram_ram_reg_56_2 : DFQD1BWP7T port map(CP => CTS_22, D => FE_PHN671_gl_ram_n_435, Q => gl_ram_ram_56(2));
  gl_ram_ram_reg_57_0 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_434, Q => gl_ram_ram_57(0));
  gl_ram_ram_reg_57_1 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_432, Q => gl_ram_ram_57(1));
  gl_ram_ram_reg_57_2 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_431, Q => gl_ram_ram_57(2));
  gl_ram_ram_reg_58_0 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_429, Q => gl_ram_ram_58(0));
  gl_ram_ram_reg_58_1 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_427, Q => FE_PHN664_gl_ram_ram_58_1);
  gl_ram_ram_reg_58_2 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_426, Q => gl_ram_ram_58(2));
  gl_ram_ram_reg_59_0 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_425, Q => gl_ram_ram_59(0));
  gl_ram_ram_reg_59_1 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_423, Q => gl_ram_ram_59(1));
  gl_ram_ram_reg_59_2 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_422, Q => FE_PHN660_gl_ram_ram_59_2);
  gl_ram_ram_reg_60_0 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_420, Q => gl_ram_ram_60(0));
  gl_ram_ram_reg_60_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_419, Q => gl_ram_ram_60(1));
  gl_ram_ram_reg_60_2 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_417, Q => gl_ram_ram_60(2));
  gl_ram_ram_reg_61_0 : DFQD1BWP7T port map(CP => CTS_22, D => gl_ram_n_416, Q => gl_ram_ram_61(0));
  gl_ram_ram_reg_61_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_414, Q => gl_ram_ram_61(1));
  gl_ram_ram_reg_61_2 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_413, Q => gl_ram_ram_61(2));
  gl_ram_ram_reg_62_0 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_411, Q => gl_ram_ram_62(0));
  gl_ram_ram_reg_62_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_409, Q => gl_ram_ram_62(1));
  gl_ram_ram_reg_62_2 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_408, Q => gl_ram_ram_62(2));
  gl_ram_ram_reg_63_0 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_407, Q => gl_ram_ram_63(0));
  gl_ram_ram_reg_63_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_405, Q => gl_ram_ram_63(1));
  gl_ram_ram_reg_63_2 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_404, Q => gl_ram_ram_63(2));
  gl_ram_ram_reg_64_0 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_295, Q => gl_ram_ram_64(0));
  gl_ram_ram_reg_64_1 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_310, Q => gl_ram_ram_64(1));
  gl_ram_ram_reg_64_2 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_293, Q => gl_ram_ram_64(2));
  gl_ram_ram_reg_65_0 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_292, Q => gl_ram_ram_65(0));
  gl_ram_ram_reg_65_1 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_291, Q => gl_ram_ram_65(1));
  gl_ram_ram_reg_65_2 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_290, Q => gl_ram_ram_65(2));
  gl_ram_ram_reg_66_0 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_289, Q => gl_ram_ram_66(0));
  gl_ram_ram_reg_66_1 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_288, Q => gl_ram_ram_66(1));
  gl_ram_ram_reg_66_2 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_287, Q => gl_ram_ram_66(2));
  gl_ram_ram_reg_67_0 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_286, Q => gl_ram_ram_67(0));
  gl_ram_ram_reg_67_1 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_285, Q => gl_ram_ram_67(1));
  gl_ram_ram_reg_67_2 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_284, Q => gl_ram_ram_67(2));
  gl_ram_ram_reg_68_0 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_283, Q => gl_ram_ram_68(0));
  gl_ram_ram_reg_68_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_282, Q => gl_ram_ram_68(1));
  gl_ram_ram_reg_68_2 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_281, Q => gl_ram_ram_68(2));
  gl_ram_ram_reg_69_0 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_280, Q => gl_ram_ram_69(0));
  gl_ram_ram_reg_69_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_294, Q => gl_ram_ram_69(1));
  gl_ram_ram_reg_69_2 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_309, Q => gl_ram_ram_69(2));
  gl_ram_ram_reg_70_0 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_277, Q => gl_ram_ram_70(0));
  gl_ram_ram_reg_70_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_276, Q => gl_ram_ram_70(1));
  gl_ram_ram_reg_70_2 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_275, Q => gl_ram_ram_70(2));
  gl_ram_ram_reg_71_0 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_274, Q => gl_ram_ram_71(0));
  gl_ram_ram_reg_71_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_273, Q => gl_ram_ram_71(1));
  gl_ram_ram_reg_71_2 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_272, Q => gl_ram_ram_71(2));
  gl_ram_ram_reg_72_0 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_271, Q => gl_ram_ram_72(0));
  gl_ram_ram_reg_72_1 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_270, Q => gl_ram_ram_72(1));
  gl_ram_ram_reg_72_2 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_269, Q => gl_ram_ram_72(2));
  gl_ram_ram_reg_73_0 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_268, Q => gl_ram_ram_73(0));
  gl_ram_ram_reg_73_1 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_267, Q => gl_ram_ram_73(1));
  gl_ram_ram_reg_73_2 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_266, Q => gl_ram_ram_73(2));
  gl_ram_ram_reg_74_0 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_265, Q => gl_ram_ram_74(0));
  gl_ram_ram_reg_74_1 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_264, Q => gl_ram_ram_74(1));
  gl_ram_ram_reg_74_2 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_263, Q => gl_ram_ram_74(2));
  gl_ram_ram_reg_75_0 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_262, Q => FE_PHN661_gl_ram_ram_75_0);
  gl_ram_ram_reg_75_1 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_261, Q => gl_ram_ram_75(1));
  gl_ram_ram_reg_75_2 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_260, Q => gl_ram_ram_75(2));
  gl_ram_ram_reg_76_0 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_259, Q => gl_ram_ram_76(0));
  gl_ram_ram_reg_76_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_258, Q => gl_ram_ram_76(1));
  gl_ram_ram_reg_76_2 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_257, Q => gl_ram_ram_76(2));
  gl_ram_ram_reg_77_0 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_256, Q => gl_ram_ram_77(0));
  gl_ram_ram_reg_77_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_255, Q => gl_ram_ram_77(1));
  gl_ram_ram_reg_77_2 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_254, Q => gl_ram_ram_77(2));
  gl_ram_ram_reg_78_0 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_253, Q => gl_ram_ram_78(0));
  gl_ram_ram_reg_78_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_252, Q => gl_ram_ram_78(1));
  gl_ram_ram_reg_78_2 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_251, Q => gl_ram_ram_78(2));
  gl_ram_ram_reg_79_0 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_250, Q => gl_ram_ram_79(0));
  gl_ram_ram_reg_79_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_249, Q => gl_ram_ram_79(1));
  gl_ram_ram_reg_79_2 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_248, Q => gl_ram_ram_79(2));
  gl_ram_ram_reg_80_0 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_378, Q => gl_ram_ram_80(0));
  gl_ram_ram_reg_80_1 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_376, Q => gl_ram_ram_80(1));
  gl_ram_ram_reg_80_2 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_375, Q => gl_ram_ram_80(2));
  gl_ram_ram_reg_81_0 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_374, Q => gl_ram_ram_81(0));
  gl_ram_ram_reg_81_1 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_372, Q => gl_ram_ram_81(1));
  gl_ram_ram_reg_81_2 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_371, Q => gl_ram_ram_81(2));
  gl_ram_ram_reg_82_0 : DFQD1BWP7T port map(CP => CTS_20, D => gl_ram_n_369, Q => gl_ram_ram_82(0));
  gl_ram_ram_reg_82_1 : DFQD1BWP7T port map(CP => CTS_20, D => gl_ram_n_368, Q => gl_ram_ram_82(1));
  gl_ram_ram_reg_82_2 : DFQD1BWP7T port map(CP => CTS_20, D => gl_ram_n_366, Q => gl_ram_ram_82(2));
  gl_ram_ram_reg_83_0 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_365, Q => gl_ram_ram_83(0));
  gl_ram_ram_reg_83_1 : DFQD1BWP7T port map(CP => CTS_20, D => gl_ram_n_363, Q => gl_ram_ram_83(1));
  gl_ram_ram_reg_83_2 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_362, Q => gl_ram_ram_83(2));
  gl_ram_ram_reg_84_0 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_360, Q => gl_ram_ram_84(0));
  gl_ram_ram_reg_84_1 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_359, Q => gl_ram_ram_84(1));
  gl_ram_ram_reg_84_2 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_357, Q => gl_ram_ram_84(2));
  gl_ram_ram_reg_85_0 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_355, Q => gl_ram_ram_85(0));
  gl_ram_ram_reg_85_1 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_353, Q => gl_ram_ram_85(1));
  gl_ram_ram_reg_85_2 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_352, Q => gl_ram_ram_85(2));
  gl_ram_ram_reg_86_0 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_350, Q => gl_ram_ram_86(0));
  gl_ram_ram_reg_86_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_348, Q => gl_ram_ram_86(1));
  gl_ram_ram_reg_86_2 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_346, Q => gl_ram_ram_86(2));
  gl_ram_ram_reg_87_0 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_345, Q => gl_ram_ram_87(0));
  gl_ram_ram_reg_87_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_343, Q => gl_ram_ram_87(1));
  gl_ram_ram_reg_87_2 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_342, Q => gl_ram_ram_87(2));
  gl_ram_ram_reg_88_0 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_341, Q => gl_ram_ram_88(0));
  gl_ram_ram_reg_88_1 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_339, Q => gl_ram_ram_88(1));
  gl_ram_ram_reg_88_2 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_337, Q => gl_ram_ram_88(2));
  gl_ram_ram_reg_89_0 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_336, Q => gl_ram_ram_89(0));
  gl_ram_ram_reg_89_1 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_334, Q => gl_ram_ram_89(1));
  gl_ram_ram_reg_89_2 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_333, Q => gl_ram_ram_89(2));
  gl_ram_ram_reg_90_0 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_331, Q => gl_ram_ram_90(0));
  gl_ram_ram_reg_90_1 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_329, Q => gl_ram_ram_90(1));
  gl_ram_ram_reg_90_2 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_327, Q => gl_ram_ram_90(2));
  gl_ram_ram_reg_91_0 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_326, Q => gl_ram_ram_91(0));
  gl_ram_ram_reg_91_1 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_324, Q => gl_ram_ram_91(1));
  gl_ram_ram_reg_91_2 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_322, Q => gl_ram_ram_91(2));
  gl_ram_ram_reg_92_0 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_320, Q => gl_ram_ram_92(0));
  gl_ram_ram_reg_92_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_319, Q => gl_ram_ram_92(1));
  gl_ram_ram_reg_92_2 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_317, Q => gl_ram_ram_92(2));
  gl_ram_ram_reg_93_0 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_316, Q => gl_ram_ram_93(0));
  gl_ram_ram_reg_93_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_314, Q => gl_ram_ram_93(1));
  gl_ram_ram_reg_93_2 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_550, Q => gl_ram_ram_93(2));
  gl_ram_ram_reg_94_0 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_549, Q => gl_ram_ram_94(0));
  gl_ram_ram_reg_94_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_547, Q => gl_ram_ram_94(1));
  gl_ram_ram_reg_94_2 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_545, Q => gl_ram_ram_94(2));
  gl_ram_ram_reg_95_0 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_544, Q => gl_ram_ram_95(0));
  gl_ram_ram_reg_95_1 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_542, Q => gl_ram_ram_95(1));
  gl_ram_ram_reg_95_2 : DFQD1BWP7T port map(CP => CTS_23, D => gl_ram_n_541, Q => gl_ram_ram_95(2));
  gl_ram_ram_reg_96_0 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_307, Q => gl_ram_ram_96(0));
  gl_ram_ram_reg_96_1 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_306, Q => gl_ram_ram_96(1));
  gl_ram_ram_reg_96_2 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_305, Q => gl_ram_ram_96(2));
  gl_ram_ram_reg_97_0 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_304, Q => gl_ram_ram_97(0));
  gl_ram_ram_reg_97_1 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_303, Q => gl_ram_ram_97(1));
  gl_ram_ram_reg_97_2 : DFQD1BWP7T port map(CP => CTS_21, D => gl_ram_n_302, Q => gl_ram_ram_97(2));
  gl_ram_ram_reg_98_0 : DFQD1BWP7T port map(CP => CTS_20, D => gl_ram_n_301, Q => gl_ram_ram_98(0));
  gl_ram_ram_reg_98_1 : DFQD1BWP7T port map(CP => CTS_20, D => gl_ram_n_300, Q => gl_ram_ram_98(1));
  gl_ram_ram_reg_98_2 : DFQD1BWP7T port map(CP => CTS_20, D => gl_ram_n_299, Q => gl_ram_ram_98(2));
  gl_ram_ram_reg_99_0 : DFQD1BWP7T port map(CP => CTS_20, D => gl_ram_n_298, Q => gl_ram_ram_99(0));
  gl_ram_ram_reg_99_1 : DFQD1BWP7T port map(CP => CTS_20, D => gl_ram_n_297, Q => gl_ram_ram_99(1));
  gl_ram_ram_reg_99_2 : DFQD1BWP7T port map(CP => CTS_20, D => gl_ram_n_296, Q => gl_ram_ram_99(2));
  gl_ram_x_grid_reg_0 : DFQD1BWP7T port map(CP => CTS_19, D => FE_PHN359_gl_ram_n_77, Q => gl_ram_x_grid(0));
  gl_ram_y_grid_reg_1 : DFQD1BWP7T port map(CP => CTS_19, D => FE_PHN370_gl_ram_n_243, Q => gl_ram_y_grid(1));
  gl_ram_g27157 : OAI211D1BWP7T port map(A1 => gl_ram_y_grid(3), A2 => gl_ram_n_140, B => gl_ram_n_565, C => gl_ram_n_555, ZN => gl_ram_n_568);
  gl_ram_g27158 : OAI31D0BWP7T port map(A1 => gl_ram_y_grid(2), A2 => gl_ram_n_4, A3 => gl_ram_n_186, B => gl_ram_n_566, ZN => FE_PHN381_gl_ram_n_567);
  gl_ram_g27159 : AOI221D0BWP7T port map(A1 => gl_ram_n_311, A2 => gl_ram_y_grid(2), B1 => gl_ram_ram_position(5), B2 => gl_ram_n_16, C => gl_ram_n_561, ZN => gl_ram_n_566);
  gl_ram_g27161 : AOI21D0BWP7T port map(A1 => gl_ram_n_232, A2 => gl_ram_n_144, B => gl_ram_n_562, ZN => gl_ram_n_565);
  gl_ram_g27163 : OR2D1BWP7T port map(A1 => gl_ram_n_559, A2 => gl_ram_n_187, Z => gl_ram_n_564);
  gl_ram_g27164 : AO221D0BWP7T port map(A1 => gl_ram_n_313, A2 => gl_ram_n_48, B1 => gl_ram_ram_position(3), B2 => gl_ram_n_16, C => gl_ram_n_560, Z => gl_ram_n_563);
  gl_ram_g27165 : OAI211D1BWP7T port map(A1 => gl_ram_n_15, A2 => gl_ram_n_0, B => gl_ram_n_558, C => gl_ram_n_312, ZN => gl_ram_n_562);
  gl_ram_g27166 : OAI22D0BWP7T port map(A1 => gl_ram_n_557, A2 => gl_ram_n_1, B1 => gl_ram_n_278, B2 => gl_ram_y_grid(2), ZN => gl_ram_n_561);
  gl_ram_g27167 : AOI31D0BWP7T port map(A1 => gl_ram_n_245, A2 => gl_ram_n_242, A3 => gl_ram_n_137, B => gl_ram_n_48, ZN => gl_ram_n_560);
  gl_ram_g27168 : OAI31D0BWP7T port map(A1 => gl_ram_x_grid(3), A2 => gl_ram_y_grid(0), A3 => gl_ram_n_231, B => gl_ram_n_556, ZN => gl_ram_n_559);
  gl_ram_g27291 : OAI222D0BWP7T port map(A1 => gl_ram_n_244, A2 => gl_ram_n_236, B1 => gl_ram_n_4, B2 => gl_ram_n_46, C1 => gl_ram_y_grid(3), C2 => gl_ram_n_18, ZN => gl_ram_n_558);
  gl_ram_g27292 : AOI222D0BWP7T port map(A1 => gl_ram_n_279, A2 => gl_ram_y_grid(3), B1 => gl_ram_n_230, B2 => gl_ram_n_6, C1 => gl_ram_n_187, C2 => gl_ram_y_grid(0), ZN => gl_ram_n_557);
  gl_ram_g27293 : MAOI22D0BWP7T port map(A1 => gl_ram_ram_position(6), A2 => gl_ram_n_16, B1 => gl_ram_n_246, B2 => gl_ram_y_grid(3), ZN => gl_ram_n_556);
  gl_ram_g27294 : AOI22D0BWP7T port map(A1 => gl_ram_n_279, A2 => gl_ram_n_79, B1 => gl_ram_n_235, B2 => gl_ram_n_240, ZN => gl_ram_n_555);
  gl_ram_g27414 : AO221D0BWP7T port map(A1 => gl_ram_n_114, A2 => gl_ram_n_111, B1 => gl_ram_n_218, B2 => FE_PHN578_gl_ram_ram_8_2, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_554);
  gl_ram_g27415 : AO221D0BWP7T port map(A1 => gl_ram_n_117, A2 => gl_ram_n_83, B1 => gl_ram_n_180, B2 => FE_PHN121_gl_ram_ram_50_0, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_553);
  gl_ram_g27416 : OAI221D0BWP7T port map(A1 => gl_ram_n_234, A2 => gl_ram_n_7, B1 => gl_ram_n_21, B2 => gl_ram_n_135, C => gl_ram_n_241, ZN => gl_ram_n_552);
  gl_ram_g27417 : AO221D0BWP7T port map(A1 => gl_ram_n_122, A2 => gl_ram_n_113, B1 => gl_ram_n_163, B2 => FE_PHN668_gl_ram_ram_1_2, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_551);
  gl_ram_g27418 : AO221D0BWP7T port map(A1 => gl_ram_n_87, A2 => gl_ram_n_81, B1 => gl_ram_n_185, B2 => FE_PHN142_gl_ram_ram_93_2, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_550);
  gl_ram_g27419 : AO221D0BWP7T port map(A1 => gl_ram_n_134, A2 => gl_ram_n_81, B1 => gl_ram_n_154, B2 => FE_PHN233_gl_ram_ram_94_0, C => gl_ram_n_16, Z => gl_ram_n_549);
  gl_ram_g27420 : AO221D0BWP7T port map(A1 => gl_ram_n_127, A2 => gl_ram_n_108, B1 => gl_ram_n_153, B2 => FE_PHN186_gl_ram_ram_30_2, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_548);
  gl_ram_g27421 : AO221D0BWP7T port map(A1 => gl_ram_n_128, A2 => gl_ram_n_81, B1 => gl_ram_n_154, B2 => FE_PHN106_gl_ram_ram_94_1, C => gl_ram_n_16, Z => gl_ram_n_547);
  gl_ram_g27422 : AO221D0BWP7T port map(A1 => gl_ram_n_126, A2 => gl_ram_n_108, B1 => gl_ram_n_147, B2 => FE_PHN172_gl_ram_ram_31_0, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_546);
  gl_ram_g27423 : AO221D0BWP7T port map(A1 => gl_ram_n_127, A2 => gl_ram_n_81, B1 => gl_ram_n_154, B2 => FE_PHN156_gl_ram_ram_94_2, C => gl_ram_n_16, Z => gl_ram_n_545);
  gl_ram_g27424 : AO221D0BWP7T port map(A1 => gl_ram_n_126, A2 => gl_ram_n_81, B1 => gl_ram_n_156, B2 => FE_PHN115_gl_ram_ram_95_0, C => gl_ram_n_16, Z => gl_ram_n_544);
  gl_ram_g27425 : AO221D0BWP7T port map(A1 => gl_ram_n_125, A2 => gl_ram_n_108, B1 => gl_ram_n_147, B2 => FE_PHN174_gl_ram_ram_31_1, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_543);
  gl_ram_g27426 : AO221D0BWP7T port map(A1 => gl_ram_n_125, A2 => gl_ram_n_81, B1 => gl_ram_n_156, B2 => FE_PHN224_gl_ram_ram_95_1, C => gl_ram_n_16, Z => gl_ram_n_542);
  gl_ram_g27427 : AO221D0BWP7T port map(A1 => gl_ram_n_129, A2 => gl_ram_n_81, B1 => gl_ram_n_156, B2 => FE_PHN259_gl_ram_ram_95_2, C => gl_ram_n_16, Z => gl_ram_n_541);
  gl_ram_g27428 : AO221D0BWP7T port map(A1 => gl_ram_n_129, A2 => gl_ram_n_108, B1 => gl_ram_n_147, B2 => FE_PHN424_gl_ram_ram_31_2, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_540);
  gl_ram_g27429 : AO221D0BWP7T port map(A1 => gl_ram_n_86, A2 => gl_ram_n_82, B1 => gl_ram_n_214, B2 => FE_PHN556_gl_ram_ram_32_0, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_539);
  gl_ram_g27430 : AO221D0BWP7T port map(A1 => gl_ram_n_117, A2 => gl_ram_n_113, B1 => gl_ram_n_166, B2 => FE_PHN569_gl_ram_ram_2_0, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_538);
  gl_ram_g27431 : AO221D0BWP7T port map(A1 => gl_ram_n_114, A2 => gl_ram_n_82, B1 => gl_ram_n_214, B2 => FE_PHN217_gl_ram_ram_32_2, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_537);
  gl_ram_g27432 : AO221D0BWP7T port map(A1 => gl_ram_n_115, A2 => gl_ram_n_82, B1 => gl_ram_n_214, B2 => FE_PHN600_gl_ram_ram_32_1, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_536);
  gl_ram_g27433 : AO221D0BWP7T port map(A1 => gl_ram_n_118, A2 => gl_ram_n_82, B1 => gl_ram_n_169, B2 => FE_PHN585_gl_ram_ram_33_0, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_535);
  gl_ram_g27434 : AO221D0BWP7T port map(A1 => gl_ram_n_120, A2 => gl_ram_n_82, B1 => gl_ram_n_169, B2 => FE_PHN427_gl_ram_ram_33_1, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_534);
  gl_ram_g27435 : AO221D0BWP7T port map(A1 => gl_ram_n_120, A2 => gl_ram_n_113, B1 => gl_ram_n_163, B2 => FE_PHN194_gl_ram_ram_1_1, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_533);
  gl_ram_g27436 : AO221D0BWP7T port map(A1 => gl_ram_n_116, A2 => gl_ram_n_113, B1 => gl_ram_n_166, B2 => FE_PHN203_gl_ram_ram_2_1, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_532);
  gl_ram_g27437 : AO221D0BWP7T port map(A1 => gl_ram_n_122, A2 => gl_ram_n_82, B1 => gl_ram_n_169, B2 => FE_PHN576_gl_ram_ram_33_2, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_531);
  gl_ram_g27438 : AO221D0BWP7T port map(A1 => gl_ram_n_117, A2 => gl_ram_n_82, B1 => gl_ram_n_168, B2 => FE_PHN187_gl_ram_ram_34_0, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_530);
  gl_ram_g27439 : AO221D0BWP7T port map(A1 => gl_ram_n_85, A2 => gl_ram_n_113, B1 => gl_ram_n_166, B2 => FE_PHN597_gl_ram_ram_2_2, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_529);
  gl_ram_g27440 : AO221D0BWP7T port map(A1 => gl_ram_n_116, A2 => gl_ram_n_82, B1 => gl_ram_n_168, B2 => FE_PHN571_gl_ram_ram_34_1, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_528);
  gl_ram_g27441 : AO221D0BWP7T port map(A1 => gl_ram_n_85, A2 => gl_ram_n_82, B1 => gl_ram_n_168, B2 => FE_PHN239_gl_ram_ram_34_2, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_527);
  gl_ram_g27442 : AO221D0BWP7T port map(A1 => gl_ram_n_119, A2 => gl_ram_n_113, B1 => gl_ram_n_162, B2 => FE_PHN562_gl_ram_ram_3_0, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_526);
  gl_ram_g27443 : AO221D0BWP7T port map(A1 => gl_ram_n_119, A2 => gl_ram_n_82, B1 => gl_ram_n_167, B2 => FE_PHN670_gl_ram_ram_35_0, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_525);
  gl_ram_g27444 : AO221D0BWP7T port map(A1 => gl_ram_n_123, A2 => gl_ram_n_82, B1 => gl_ram_n_167, B2 => FE_PHN169_gl_ram_ram_35_1, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_524);
  gl_ram_g27445 : AO221D0BWP7T port map(A1 => gl_ram_n_121, A2 => gl_ram_n_82, B1 => gl_ram_n_167, B2 => FE_PHN592_gl_ram_ram_35_2, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_523);
  gl_ram_g27446 : AO221D0BWP7T port map(A1 => gl_ram_n_133, A2 => gl_ram_n_82, B1 => gl_ram_n_204, B2 => FE_PHN274_gl_ram_ram_36_0, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_522);
  gl_ram_g27447 : AO221D0BWP7T port map(A1 => gl_ram_n_132, A2 => gl_ram_n_82, B1 => gl_ram_n_204, B2 => FE_PHN285_gl_ram_ram_36_1, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_521);
  gl_ram_g27448 : AO221D0BWP7T port map(A1 => gl_ram_n_131, A2 => gl_ram_n_82, B1 => gl_ram_n_204, B2 => FE_PHN428_gl_ram_ram_36_2, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_520);
  gl_ram_g27449 : AO221D0BWP7T port map(A1 => gl_ram_n_123, A2 => gl_ram_n_113, B1 => gl_ram_n_162, B2 => FE_PHN171_gl_ram_ram_3_1, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_519);
  gl_ram_g27450 : AO221D0BWP7T port map(A1 => gl_ram_n_124, A2 => gl_ram_n_82, B1 => gl_ram_n_208, B2 => FE_PHN309_gl_ram_ram_37_0, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_518);
  gl_ram_g27451 : AO221D0BWP7T port map(A1 => gl_ram_n_121, A2 => gl_ram_n_113, B1 => gl_ram_n_162, B2 => FE_PHN567_gl_ram_ram_3_2, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_517);
  gl_ram_g27452 : AO221D0BWP7T port map(A1 => gl_ram_n_130, A2 => gl_ram_n_82, B1 => gl_ram_n_208, B2 => FE_PHN127_gl_ram_ram_37_1, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_516);
  gl_ram_g27453 : AO221D0BWP7T port map(A1 => gl_ram_n_87, A2 => gl_ram_n_82, B1 => gl_ram_n_208, B2 => FE_PHN662_gl_ram_ram_37_2, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_515);
  gl_ram_g27454 : AO221D0BWP7T port map(A1 => gl_ram_n_133, A2 => gl_ram_n_113, B1 => gl_ram_n_205, B2 => FE_PHN507_gl_ram_ram_4_0, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_514);
  gl_ram_g27455 : AO221D0BWP7T port map(A1 => gl_ram_n_134, A2 => gl_ram_n_82, B1 => gl_ram_n_207, B2 => FE_PHN146_gl_ram_ram_38_0, C => gl_ram_n_16, Z => gl_ram_n_513);
  gl_ram_g27456 : AO221D0BWP7T port map(A1 => gl_ram_n_128, A2 => gl_ram_n_82, B1 => gl_ram_n_207, B2 => FE_PHN288_gl_ram_ram_38_1, C => gl_ram_n_16, Z => gl_ram_n_512);
  gl_ram_g27457 : AO221D0BWP7T port map(A1 => gl_ram_n_127, A2 => gl_ram_n_82, B1 => gl_ram_n_207, B2 => FE_PHN202_gl_ram_ram_38_2, C => gl_ram_n_16, Z => gl_ram_n_511);
  gl_ram_g27458 : AO221D0BWP7T port map(A1 => gl_ram_n_126, A2 => gl_ram_n_82, B1 => gl_ram_n_209, B2 => FE_PHN293_gl_ram_ram_39_0, C => gl_ram_n_16, Z => gl_ram_n_510);
  gl_ram_g27459 : AO221D0BWP7T port map(A1 => gl_ram_n_132, A2 => gl_ram_n_113, B1 => gl_ram_n_205, B2 => FE_PHN243_gl_ram_ram_4_1, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_509);
  gl_ram_g27460 : AO221D0BWP7T port map(A1 => gl_ram_n_131, A2 => gl_ram_n_113, B1 => gl_ram_n_205, B2 => FE_PHN94_gl_ram_ram_4_2, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_508);
  gl_ram_g27461 : AO221D0BWP7T port map(A1 => gl_ram_n_125, A2 => gl_ram_n_82, B1 => gl_ram_n_209, B2 => FE_PHN180_gl_ram_ram_39_1, C => gl_ram_n_16, Z => gl_ram_n_507);
  gl_ram_g27462 : AO221D0BWP7T port map(A1 => gl_ram_n_129, A2 => gl_ram_n_82, B1 => gl_ram_n_209, B2 => FE_PHN306_gl_ram_ram_39_2, C => gl_ram_n_16, Z => gl_ram_n_506);
  gl_ram_g27463 : AO221D0BWP7T port map(A1 => gl_ram_n_86, A2 => gl_ram_n_110, B1 => gl_ram_n_215, B2 => FE_PHN554_gl_ram_ram_40_0, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_505);
  gl_ram_g27464 : AO221D0BWP7T port map(A1 => gl_ram_n_115, A2 => gl_ram_n_110, B1 => gl_ram_n_215, B2 => FE_PHN527_gl_ram_ram_40_1, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_504);
  gl_ram_g27465 : AO221D0BWP7T port map(A1 => gl_ram_n_124, A2 => gl_ram_n_113, B1 => gl_ram_n_175, B2 => FE_PHN442_gl_ram_ram_5_0, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_503);
  gl_ram_g27466 : AO221D0BWP7T port map(A1 => gl_ram_n_114, A2 => gl_ram_n_110, B1 => gl_ram_n_215, B2 => FE_PHN163_gl_ram_ram_40_2, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_502);
  gl_ram_g27467 : AO221D0BWP7T port map(A1 => gl_ram_n_118, A2 => gl_ram_n_110, B1 => gl_ram_n_157, B2 => FE_PHN582_gl_ram_ram_41_0, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_501);
  gl_ram_g27468 : AO221D0BWP7T port map(A1 => gl_ram_n_120, A2 => gl_ram_n_110, B1 => gl_ram_n_157, B2 => FE_PHN222_gl_ram_ram_41_1, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_500);
  gl_ram_g27469 : AO221D0BWP7T port map(A1 => gl_ram_n_122, A2 => gl_ram_n_110, B1 => gl_ram_n_157, B2 => FE_PHN411_gl_ram_ram_41_2, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_499);
  gl_ram_g27470 : AO221D0BWP7T port map(A1 => gl_ram_n_130, A2 => gl_ram_n_113, B1 => gl_ram_n_175, B2 => FE_PHN492_gl_ram_ram_5_1, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_498);
  gl_ram_g27471 : AO221D0BWP7T port map(A1 => gl_ram_n_117, A2 => gl_ram_n_110, B1 => gl_ram_n_149, B2 => FE_PHN167_gl_ram_ram_42_0, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_497);
  gl_ram_g27472 : AO221D0BWP7T port map(A1 => gl_ram_n_116, A2 => gl_ram_n_110, B1 => gl_ram_n_149, B2 => gl_ram_ram_42(1), C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_496);
  gl_ram_g27473 : AO221D0BWP7T port map(A1 => gl_ram_n_85, A2 => gl_ram_n_110, B1 => gl_ram_n_149, B2 => gl_ram_ram_42(2), C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_495);
  gl_ram_g27474 : AO221D0BWP7T port map(A1 => gl_ram_n_119, A2 => gl_ram_n_110, B1 => gl_ram_n_150, B2 => FE_PHN559_gl_ram_ram_43_0, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_494);
  gl_ram_g27475 : AO221D0BWP7T port map(A1 => gl_ram_n_134, A2 => gl_ram_n_113, B1 => gl_ram_n_174, B2 => FE_PHN269_gl_ram_ram_6_0, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_493);
  gl_ram_g27476 : AO221D0BWP7T port map(A1 => gl_ram_n_123, A2 => gl_ram_n_110, B1 => gl_ram_n_150, B2 => FE_PHN525_gl_ram_ram_43_1, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_492);
  gl_ram_g27477 : AO221D0BWP7T port map(A1 => gl_ram_n_87, A2 => gl_ram_n_113, B1 => gl_ram_n_175, B2 => FE_PHN102_gl_ram_ram_5_2, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_491);
  gl_ram_g27478 : AO221D0BWP7T port map(A1 => gl_ram_n_121, A2 => gl_ram_n_110, B1 => gl_ram_n_150, B2 => FE_PHN564_gl_ram_ram_43_2, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_490);
  gl_ram_g27479 : AO221D0BWP7T port map(A1 => gl_ram_n_133, A2 => gl_ram_n_110, B1 => gl_ram_n_203, B2 => gl_ram_ram_44(0), C => FE_OFN38_gl_ram_n_16, Z => FE_PHN579_gl_ram_n_489);
  gl_ram_g27480 : AO221D0BWP7T port map(A1 => gl_ram_n_132, A2 => gl_ram_n_110, B1 => gl_ram_n_203, B2 => FE_PHN111_gl_ram_ram_44_1, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_488);
  gl_ram_g27481 : AO221D0BWP7T port map(A1 => gl_ram_n_131, A2 => gl_ram_n_110, B1 => gl_ram_n_203, B2 => FE_PHN225_gl_ram_ram_44_2, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_487);
  gl_ram_g27482 : AO221D0BWP7T port map(A1 => gl_ram_n_128, A2 => gl_ram_n_113, B1 => gl_ram_n_174, B2 => FE_PHN268_gl_ram_ram_6_1, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_486);
  gl_ram_g27483 : AO221D0BWP7T port map(A1 => gl_ram_n_127, A2 => gl_ram_n_113, B1 => gl_ram_n_174, B2 => FE_PHN263_gl_ram_ram_6_2, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_485);
  gl_ram_g27484 : AO221D0BWP7T port map(A1 => gl_ram_n_124, A2 => gl_ram_n_110, B1 => gl_ram_n_210, B2 => FE_PHN120_gl_ram_ram_45_0, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_484);
  gl_ram_g27485 : AO221D0BWP7T port map(A1 => gl_ram_n_130, A2 => gl_ram_n_110, B1 => gl_ram_n_210, B2 => FE_PHN260_gl_ram_ram_45_1, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_483);
  gl_ram_g27486 : AO221D0BWP7T port map(A1 => gl_ram_n_87, A2 => gl_ram_n_110, B1 => gl_ram_n_210, B2 => FE_PHN145_gl_ram_ram_45_2, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_482);
  gl_ram_g27487 : AO221D0BWP7T port map(A1 => gl_ram_n_126, A2 => gl_ram_n_113, B1 => gl_ram_n_178, B2 => FE_PHN195_gl_ram_ram_7_0, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_481);
  gl_ram_g27488 : AO221D0BWP7T port map(A1 => gl_ram_n_134, A2 => gl_ram_n_110, B1 => gl_ram_n_211, B2 => FE_PHN138_gl_ram_ram_46_0, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_480);
  gl_ram_g27489 : AO221D0BWP7T port map(A1 => gl_ram_n_125, A2 => gl_ram_n_113, B1 => gl_ram_n_178, B2 => FE_PHN173_gl_ram_ram_7_1, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_479);
  gl_ram_g27490 : AO221D0BWP7T port map(A1 => gl_ram_n_128, A2 => gl_ram_n_110, B1 => gl_ram_n_211, B2 => FE_PHN289_gl_ram_ram_46_1, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_478);
  gl_ram_g27491 : AO221D0BWP7T port map(A1 => gl_ram_n_127, A2 => gl_ram_n_110, B1 => gl_ram_n_211, B2 => FE_PHN449_gl_ram_ram_46_2, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_477);
  gl_ram_g27492 : AO221D0BWP7T port map(A1 => gl_ram_n_126, A2 => gl_ram_n_110, B1 => gl_ram_n_212, B2 => FE_PHN272_gl_ram_ram_47_0, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_476);
  gl_ram_g27493 : AO221D0BWP7T port map(A1 => gl_ram_n_125, A2 => gl_ram_n_110, B1 => gl_ram_n_212, B2 => FE_PHN231_gl_ram_ram_47_1, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_475);
  gl_ram_g27494 : AO221D0BWP7T port map(A1 => gl_ram_n_129, A2 => gl_ram_n_113, B1 => gl_ram_n_178, B2 => FE_PHN95_gl_ram_ram_7_2, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_474);
  gl_ram_g27495 : AO221D0BWP7T port map(A1 => gl_ram_n_129, A2 => gl_ram_n_110, B1 => gl_ram_n_212, B2 => FE_PHN206_gl_ram_ram_47_2, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_473);
  gl_ram_g27496 : AO221D0BWP7T port map(A1 => gl_ram_n_86, A2 => gl_ram_n_83, B1 => gl_ram_n_223, B2 => FE_PHN165_gl_ram_ram_48_0, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_472);
  gl_ram_g27497 : AO221D0BWP7T port map(A1 => gl_ram_n_115, A2 => gl_ram_n_83, B1 => gl_ram_n_223, B2 => FE_PHN637_gl_ram_ram_48_1, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_471);
  gl_ram_g27498 : AO221D0BWP7T port map(A1 => gl_ram_n_86, A2 => gl_ram_n_111, B1 => gl_ram_n_218, B2 => FE_PHN575_gl_ram_ram_8_0, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_470);
  gl_ram_g27499 : AO221D0BWP7T port map(A1 => gl_ram_n_114, A2 => gl_ram_n_83, B1 => gl_ram_n_223, B2 => FE_PHN533_gl_ram_ram_48_2, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_469);
  gl_ram_g27500 : AO221D0BWP7T port map(A1 => gl_ram_n_118, A2 => gl_ram_n_83, B1 => gl_ram_n_181, B2 => FE_PHN213_gl_ram_ram_49_0, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_468);
  gl_ram_g27501 : AO221D0BWP7T port map(A1 => gl_ram_n_115, A2 => gl_ram_n_111, B1 => gl_ram_n_218, B2 => FE_PHN572_gl_ram_ram_8_1, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_467);
  gl_ram_g27502 : AO221D0BWP7T port map(A1 => gl_ram_n_120, A2 => gl_ram_n_83, B1 => gl_ram_n_181, B2 => FE_PHN227_gl_ram_ram_49_1, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_466);
  gl_ram_g27503 : AO221D0BWP7T port map(A1 => gl_ram_n_122, A2 => gl_ram_n_83, B1 => gl_ram_n_181, B2 => FE_PHN208_gl_ram_ram_49_2, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_465);
  gl_ram_g27504 : AO221D0BWP7T port map(A1 => gl_ram_n_116, A2 => gl_ram_n_83, B1 => gl_ram_n_180, B2 => FE_PHN633_gl_ram_ram_50_1, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_464);
  gl_ram_g27567 : AO221D0BWP7T port map(A1 => gl_ram_n_85, A2 => gl_ram_n_83, B1 => gl_ram_n_180, B2 => FE_PHN634_gl_ram_ram_50_2, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_463);
  gl_ram_g27568 : AO221D0BWP7T port map(A1 => gl_ram_n_119, A2 => gl_ram_n_83, B1 => gl_ram_n_179, B2 => FE_PHN179_gl_ram_ram_51_0, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_462);
  gl_ram_g27569 : AO221D0BWP7T port map(A1 => gl_ram_n_120, A2 => gl_ram_n_111, B1 => gl_ram_n_164, B2 => FE_PHN149_gl_ram_ram_9_1, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_461);
  gl_ram_g27570 : AO221D0BWP7T port map(A1 => gl_ram_n_123, A2 => gl_ram_n_83, B1 => gl_ram_n_179, B2 => FE_PHN122_gl_ram_ram_51_1, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_460);
  gl_ram_g27571 : AO221D0BWP7T port map(A1 => gl_ram_n_121, A2 => gl_ram_n_83, B1 => gl_ram_n_179, B2 => FE_PHN586_gl_ram_ram_51_2, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_459);
  gl_ram_g27572 : AO221D0BWP7T port map(A1 => gl_ram_n_118, A2 => gl_ram_n_111, B1 => gl_ram_n_164, B2 => FE_PHN565_gl_ram_ram_9_0, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_458);
  gl_ram_g27573 : AO221D0BWP7T port map(A1 => gl_ram_n_122, A2 => gl_ram_n_111, B1 => gl_ram_n_164, B2 => FE_PHN648_gl_ram_ram_9_2, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_457);
  gl_ram_g27574 : AO221D0BWP7T port map(A1 => gl_ram_n_133, A2 => gl_ram_n_83, B1 => gl_ram_n_216, B2 => FE_PHN178_gl_ram_ram_52_0, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_456);
  gl_ram_g27575 : AO221D0BWP7T port map(A1 => gl_ram_n_132, A2 => gl_ram_n_83, B1 => gl_ram_n_216, B2 => FE_PHN133_gl_ram_ram_52_1, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_455);
  gl_ram_g27576 : AO221D0BWP7T port map(A1 => gl_ram_n_117, A2 => gl_ram_n_111, B1 => gl_ram_n_165, B2 => FE_PHN438_gl_ram_ram_10_0, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_454);
  gl_ram_g27577 : AO221D0BWP7T port map(A1 => gl_ram_n_131, A2 => gl_ram_n_83, B1 => gl_ram_n_216, B2 => FE_PHN278_gl_ram_ram_52_2, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_453);
  gl_ram_g27578 : AO221D0BWP7T port map(A1 => gl_ram_n_124, A2 => gl_ram_n_83, B1 => gl_ram_n_173, B2 => FE_PHN290_gl_ram_ram_53_0, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_452);
  gl_ram_g27579 : AO221D0BWP7T port map(A1 => gl_ram_n_116, A2 => gl_ram_n_111, B1 => gl_ram_n_165, B2 => FE_PHN160_gl_ram_ram_10_1, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_451);
  gl_ram_g27580 : AO221D0BWP7T port map(A1 => gl_ram_n_130, A2 => gl_ram_n_83, B1 => gl_ram_n_173, B2 => FE_PHN283_gl_ram_ram_53_1, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_450);
  gl_ram_g27581 : AO221D0BWP7T port map(A1 => gl_ram_n_87, A2 => gl_ram_n_83, B1 => gl_ram_n_173, B2 => FE_PHN117_gl_ram_ram_53_2, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_449);
  gl_ram_g27582 : AO221D0BWP7T port map(A1 => gl_ram_n_85, A2 => gl_ram_n_111, B1 => gl_ram_n_165, B2 => FE_PHN166_gl_ram_ram_10_2, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_448);
  gl_ram_g27583 : AO221D0BWP7T port map(A1 => gl_ram_n_134, A2 => gl_ram_n_83, B1 => gl_ram_n_172, B2 => FE_PHN100_gl_ram_ram_54_0, C => gl_ram_n_16, Z => gl_ram_n_447);
  gl_ram_g27584 : AO221D0BWP7T port map(A1 => gl_ram_n_128, A2 => gl_ram_n_83, B1 => gl_ram_n_172, B2 => FE_PHN261_gl_ram_ram_54_1, C => gl_ram_n_16, Z => gl_ram_n_446);
  gl_ram_g27585 : AO221D0BWP7T port map(A1 => gl_ram_n_119, A2 => gl_ram_n_111, B1 => gl_ram_n_161, B2 => FE_PHN532_gl_ram_ram_11_0, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_445);
  gl_ram_g27586 : AO221D0BWP7T port map(A1 => gl_ram_n_127, A2 => gl_ram_n_83, B1 => gl_ram_n_172, B2 => FE_PHN198_gl_ram_ram_54_2, C => gl_ram_n_16, Z => gl_ram_n_444);
  gl_ram_g27587 : AO221D0BWP7T port map(A1 => gl_ram_n_126, A2 => gl_ram_n_83, B1 => gl_ram_n_176, B2 => FE_PHN249_gl_ram_ram_55_0, C => gl_ram_n_16, Z => gl_ram_n_443);
  gl_ram_g27588 : AO221D0BWP7T port map(A1 => gl_ram_n_123, A2 => gl_ram_n_111, B1 => gl_ram_n_161, B2 => FE_PHN568_gl_ram_ram_11_1, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_442);
  gl_ram_g27589 : AO221D0BWP7T port map(A1 => gl_ram_n_125, A2 => gl_ram_n_83, B1 => gl_ram_n_176, B2 => FE_PHN276_gl_ram_ram_55_1, C => gl_ram_n_16, Z => gl_ram_n_441);
  gl_ram_g27590 : AO221D0BWP7T port map(A1 => gl_ram_n_129, A2 => gl_ram_n_83, B1 => gl_ram_n_176, B2 => FE_PHN262_gl_ram_ram_55_2, C => gl_ram_n_16, Z => gl_ram_n_440);
  gl_ram_g27591 : AO221D0BWP7T port map(A1 => gl_ram_n_121, A2 => gl_ram_n_111, B1 => gl_ram_n_161, B2 => FE_PHN510_gl_ram_ram_11_2, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_439);
  gl_ram_g27592 : AO221D0BWP7T port map(A1 => gl_ram_n_86, A2 => gl_ram_n_109, B1 => gl_ram_n_213, B2 => FE_PHN148_gl_ram_ram_56_0, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_438);
  gl_ram_g27593 : AO221D0BWP7T port map(A1 => gl_ram_n_115, A2 => gl_ram_n_109, B1 => gl_ram_n_213, B2 => FE_PHN590_gl_ram_ram_56_1, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_437);
  gl_ram_g27594 : AO221D0BWP7T port map(A1 => gl_ram_n_133, A2 => gl_ram_n_111, B1 => gl_ram_n_206, B2 => FE_PHN140_gl_ram_ram_12_0, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_436);
  gl_ram_g27595 : AO221D0BWP7T port map(A1 => gl_ram_n_114, A2 => gl_ram_n_109, B1 => gl_ram_n_213, B2 => FE_PHN591_gl_ram_ram_56_2, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_435);
  gl_ram_g27596 : AO221D0BWP7T port map(A1 => gl_ram_n_118, A2 => gl_ram_n_109, B1 => gl_ram_n_158, B2 => FE_PHN211_gl_ram_ram_57_0, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_434);
  gl_ram_g27597 : AO221D0BWP7T port map(A1 => gl_ram_n_132, A2 => gl_ram_n_111, B1 => gl_ram_n_206, B2 => FE_PHN595_gl_ram_ram_12_1, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_433);
  gl_ram_g27598 : AO221D0BWP7T port map(A1 => gl_ram_n_120, A2 => gl_ram_n_109, B1 => gl_ram_n_158, B2 => FE_PHN632_gl_ram_ram_57_1, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_432);
  gl_ram_g27599 : AO221D0BWP7T port map(A1 => gl_ram_n_122, A2 => gl_ram_n_109, B1 => gl_ram_n_158, B2 => FE_PHN134_gl_ram_ram_57_2, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_431);
  gl_ram_g27600 : AO221D0BWP7T port map(A1 => gl_ram_n_131, A2 => gl_ram_n_111, B1 => gl_ram_n_206, B2 => FE_PHN644_gl_ram_ram_12_2, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_430);
  gl_ram_g27601 : AO221D0BWP7T port map(A1 => gl_ram_n_117, A2 => gl_ram_n_109, B1 => gl_ram_n_159, B2 => FE_PHN185_gl_ram_ram_58_0, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_429);
  gl_ram_g27602 : AO221D0BWP7T port map(A1 => gl_ram_n_124, A2 => gl_ram_n_111, B1 => gl_ram_n_171, B2 => FE_PHN266_gl_ram_ram_13_0, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_428);
  gl_ram_g27603 : AO221D0BWP7T port map(A1 => gl_ram_n_116, A2 => gl_ram_n_109, B1 => gl_ram_n_159, B2 => FE_PHN606_gl_ram_ram_58_1, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_427);
  gl_ram_g27604 : AO221D0BWP7T port map(A1 => gl_ram_n_85, A2 => gl_ram_n_109, B1 => gl_ram_n_159, B2 => FE_PHN247_gl_ram_ram_58_2, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_426);
  gl_ram_g27605 : AO221D0BWP7T port map(A1 => gl_ram_n_119, A2 => gl_ram_n_109, B1 => gl_ram_n_160, B2 => FE_PHN228_gl_ram_ram_59_0, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_425);
  gl_ram_g27606 : AO221D0BWP7T port map(A1 => gl_ram_n_130, A2 => gl_ram_n_111, B1 => gl_ram_n_171, B2 => FE_PHN126_gl_ram_ram_13_1, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_424);
  gl_ram_g27607 : AO221D0BWP7T port map(A1 => gl_ram_n_123, A2 => gl_ram_n_109, B1 => gl_ram_n_160, B2 => FE_PHN118_gl_ram_ram_59_1, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_423);
  gl_ram_g27608 : AO221D0BWP7T port map(A1 => gl_ram_n_121, A2 => gl_ram_n_109, B1 => gl_ram_n_160, B2 => FE_PHN485_gl_ram_ram_59_2, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_422);
  gl_ram_g27609 : AO221D0BWP7T port map(A1 => gl_ram_n_87, A2 => gl_ram_n_111, B1 => gl_ram_n_171, B2 => FE_PHN177_gl_ram_ram_13_2, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_421);
  gl_ram_g27610 : AO221D0BWP7T port map(A1 => gl_ram_n_133, A2 => gl_ram_n_109, B1 => gl_ram_n_202, B2 => FE_PHN431_gl_ram_ram_60_0, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_420);
  gl_ram_g27611 : AO221D0BWP7T port map(A1 => gl_ram_n_132, A2 => gl_ram_n_109, B1 => gl_ram_n_202, B2 => FE_PHN429_gl_ram_ram_60_1, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_419);
  gl_ram_g27612 : AO221D0BWP7T port map(A1 => gl_ram_n_134, A2 => gl_ram_n_111, B1 => gl_ram_n_170, B2 => FE_PHN292_gl_ram_ram_14_0, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_418);
  gl_ram_g27613 : AO221D0BWP7T port map(A1 => gl_ram_n_131, A2 => gl_ram_n_109, B1 => gl_ram_n_202, B2 => FE_PHN430_gl_ram_ram_60_2, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_417);
  gl_ram_g27614 : AO221D0BWP7T port map(A1 => gl_ram_n_124, A2 => gl_ram_n_109, B1 => gl_ram_n_228, B2 => FE_PHN253_gl_ram_ram_61_0, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_416);
  gl_ram_g27615 : AO221D0BWP7T port map(A1 => gl_ram_n_128, A2 => gl_ram_n_111, B1 => gl_ram_n_170, B2 => FE_PHN205_gl_ram_ram_14_1, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_415);
  gl_ram_g27616 : AO221D0BWP7T port map(A1 => gl_ram_n_130, A2 => gl_ram_n_109, B1 => gl_ram_n_228, B2 => FE_PHN439_gl_ram_ram_61_1, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_414);
  gl_ram_g27617 : AO221D0BWP7T port map(A1 => gl_ram_n_87, A2 => gl_ram_n_109, B1 => gl_ram_n_228, B2 => FE_PHN244_gl_ram_ram_61_2, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_413);
  gl_ram_g27618 : AO221D0BWP7T port map(A1 => gl_ram_n_127, A2 => gl_ram_n_111, B1 => gl_ram_n_170, B2 => FE_PHN295_gl_ram_ram_14_2, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_412);
  gl_ram_g27619 : AO221D0BWP7T port map(A1 => gl_ram_n_134, A2 => gl_ram_n_109, B1 => gl_ram_n_229, B2 => FE_PHN124_gl_ram_ram_62_0, C => gl_ram_n_16, Z => gl_ram_n_411);
  gl_ram_g27620 : AO221D0BWP7T port map(A1 => gl_ram_n_126, A2 => gl_ram_n_111, B1 => gl_ram_n_177, B2 => FE_PHN204_gl_ram_ram_15_0, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_410);
  gl_ram_g27621 : AO221D0BWP7T port map(A1 => gl_ram_n_128, A2 => gl_ram_n_109, B1 => gl_ram_n_229, B2 => FE_PHN232_gl_ram_ram_62_1, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_409);
  gl_ram_g27622 : AO221D0BWP7T port map(A1 => gl_ram_n_127, A2 => gl_ram_n_109, B1 => gl_ram_n_229, B2 => FE_PHN207_gl_ram_ram_62_2, C => gl_ram_n_16, Z => gl_ram_n_408);
  gl_ram_g27623 : AO221D0BWP7T port map(A1 => gl_ram_n_126, A2 => gl_ram_n_109, B1 => gl_ram_n_189, B2 => FE_PHN273_gl_ram_ram_63_0, C => gl_ram_n_16, Z => gl_ram_n_407);
  gl_ram_g27624 : AO221D0BWP7T port map(A1 => gl_ram_n_125, A2 => gl_ram_n_111, B1 => gl_ram_n_177, B2 => FE_PHN175_gl_ram_ram_15_1, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_406);
  gl_ram_g27625 : AO221D0BWP7T port map(A1 => gl_ram_n_125, A2 => gl_ram_n_109, B1 => gl_ram_n_189, B2 => FE_PHN277_gl_ram_ram_63_1, C => gl_ram_n_16, Z => gl_ram_n_405);
  gl_ram_g27626 : AO221D0BWP7T port map(A1 => gl_ram_n_129, A2 => gl_ram_n_109, B1 => gl_ram_n_189, B2 => FE_PHN254_gl_ram_ram_63_2, C => gl_ram_n_16, Z => gl_ram_n_404);
  gl_ram_g27627 : AO221D0BWP7T port map(A1 => gl_ram_n_129, A2 => gl_ram_n_111, B1 => gl_ram_n_177, B2 => FE_PHN267_gl_ram_ram_15_2, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_403);
  gl_ram_g27628 : AO221D0BWP7T port map(A1 => gl_ram_n_86, A2 => gl_ram_n_112, B1 => gl_ram_n_226, B2 => FE_PHN192_gl_ram_ram_16_0, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_402);
  gl_ram_g27629 : AO221D0BWP7T port map(A1 => gl_ram_n_115, A2 => gl_ram_n_112, B1 => gl_ram_n_226, B2 => FE_PHN97_gl_ram_ram_16_1, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_401);
  gl_ram_g27630 : AO221D0BWP7T port map(A1 => gl_ram_n_114, A2 => gl_ram_n_112, B1 => gl_ram_n_226, B2 => FE_PHN598_gl_ram_ram_16_2, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_400);
  gl_ram_g27631 : AO221D0BWP7T port map(A1 => gl_ram_n_118, A2 => gl_ram_n_112, B1 => gl_ram_n_198, B2 => FE_PHN131_gl_ram_ram_17_0, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_399);
  gl_ram_g27632 : AO221D0BWP7T port map(A1 => gl_ram_n_120, A2 => gl_ram_n_112, B1 => gl_ram_n_198, B2 => FE_PHN511_gl_ram_ram_17_1, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_398);
  gl_ram_g27633 : AO221D0BWP7T port map(A1 => gl_ram_n_122, A2 => gl_ram_n_112, B1 => gl_ram_n_198, B2 => FE_PHN96_gl_ram_ram_17_2, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_397);
  gl_ram_g27634 : AO221D0BWP7T port map(A1 => gl_ram_n_117, A2 => gl_ram_n_112, B1 => gl_ram_n_195, B2 => FE_PHN659_gl_ram_ram_18_0, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_396);
  gl_ram_g27635 : AO221D0BWP7T port map(A1 => gl_ram_n_116, A2 => gl_ram_n_112, B1 => gl_ram_n_195, B2 => FE_PHN136_gl_ram_ram_18_1, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_395);
  gl_ram_g27636 : AO221D0BWP7T port map(A1 => gl_ram_n_85, A2 => gl_ram_n_112, B1 => gl_ram_n_195, B2 => gl_ram_ram_18(2), C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_394);
  gl_ram_g27637 : AO221D0BWP7T port map(A1 => gl_ram_n_119, A2 => gl_ram_n_112, B1 => gl_ram_n_191, B2 => FE_PHN558_gl_ram_ram_19_0, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_393);
  gl_ram_g27638 : AO221D0BWP7T port map(A1 => gl_ram_n_123, A2 => gl_ram_n_112, B1 => gl_ram_n_191, B2 => FE_PHN476_gl_ram_ram_19_1, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_392);
  gl_ram_g27639 : AO221D0BWP7T port map(A1 => gl_ram_n_121, A2 => gl_ram_n_112, B1 => gl_ram_n_191, B2 => FE_PHN158_gl_ram_ram_19_2, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_391);
  gl_ram_g27640 : AO221D0BWP7T port map(A1 => gl_ram_n_133, A2 => gl_ram_n_112, B1 => gl_ram_n_221, B2 => FE_PHN245_gl_ram_ram_20_0, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_390);
  gl_ram_g27641 : AO221D0BWP7T port map(A1 => gl_ram_n_132, A2 => gl_ram_n_112, B1 => gl_ram_n_221, B2 => FE_PHN422_gl_ram_ram_20_1, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_389);
  gl_ram_g27642 : AO221D0BWP7T port map(A1 => gl_ram_n_131, A2 => gl_ram_n_112, B1 => gl_ram_n_221, B2 => FE_PHN450_gl_ram_ram_20_2, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_388);
  gl_ram_g27643 : AO221D0BWP7T port map(A1 => gl_ram_n_124, A2 => gl_ram_n_112, B1 => gl_ram_n_155, B2 => FE_PHN601_gl_ram_ram_21_0, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_387);
  gl_ram_g27644 : AO221D0BWP7T port map(A1 => gl_ram_n_130, A2 => gl_ram_n_112, B1 => gl_ram_n_155, B2 => FE_PHN184_gl_ram_ram_21_1, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_386);
  gl_ram_g27645 : AO221D0BWP7T port map(A1 => gl_ram_n_87, A2 => gl_ram_n_112, B1 => gl_ram_n_155, B2 => FE_PHN105_gl_ram_ram_21_2, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_385);
  gl_ram_g27646 : AO221D0BWP7T port map(A1 => gl_ram_n_134, A2 => gl_ram_n_112, B1 => gl_ram_n_151, B2 => FE_PHN265_gl_ram_ram_22_0, C => gl_ram_n_16, Z => gl_ram_n_384);
  gl_ram_g27647 : AO221D0BWP7T port map(A1 => gl_ram_n_128, A2 => gl_ram_n_112, B1 => gl_ram_n_151, B2 => FE_PHN281_gl_ram_ram_22_1, C => gl_ram_n_16, Z => gl_ram_n_383);
  gl_ram_g27648 : AO221D0BWP7T port map(A1 => gl_ram_n_127, A2 => gl_ram_n_112, B1 => gl_ram_n_151, B2 => FE_PHN183_gl_ram_ram_22_2, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_382);
  gl_ram_g27649 : AO221D0BWP7T port map(A1 => gl_ram_n_126, A2 => gl_ram_n_112, B1 => gl_ram_n_183, B2 => FE_PHN155_gl_ram_ram_23_0, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_381);
  gl_ram_g27650 : AO221D0BWP7T port map(A1 => gl_ram_n_125, A2 => gl_ram_n_112, B1 => gl_ram_n_183, B2 => FE_PHN282_gl_ram_ram_23_1, C => gl_ram_n_16, Z => gl_ram_n_380);
  gl_ram_g27651 : AO221D0BWP7T port map(A1 => gl_ram_n_129, A2 => gl_ram_n_112, B1 => gl_ram_n_183, B2 => FE_PHN287_gl_ram_ram_23_2, C => gl_ram_n_16, Z => gl_ram_n_379);
  gl_ram_g27652 : AO221D0BWP7T port map(A1 => gl_ram_n_86, A2 => gl_ram_n_84, B1 => gl_ram_n_225, B2 => FE_PHN444_gl_ram_ram_80_0, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_378);
  gl_ram_g27653 : AO221D0BWP7T port map(A1 => gl_ram_n_86, A2 => gl_ram_n_108, B1 => gl_ram_n_227, B2 => FE_PHN563_gl_ram_ram_24_0, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_377);
  gl_ram_g27654 : AO221D0BWP7T port map(A1 => gl_ram_n_115, A2 => gl_ram_n_84, B1 => gl_ram_n_225, B2 => FE_PHN132_gl_ram_ram_80_1, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_376);
  gl_ram_g27655 : AO221D0BWP7T port map(A1 => gl_ram_n_114, A2 => gl_ram_n_84, B1 => gl_ram_n_225, B2 => FE_PHN209_gl_ram_ram_80_2, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_375);
  gl_ram_g27656 : AO221D0BWP7T port map(A1 => gl_ram_n_118, A2 => gl_ram_n_84, B1 => gl_ram_n_200, B2 => FE_PHN150_gl_ram_ram_81_0, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_374);
  gl_ram_g27657 : AO221D0BWP7T port map(A1 => gl_ram_n_115, A2 => gl_ram_n_108, B1 => gl_ram_n_227, B2 => FE_PHN557_gl_ram_ram_24_1, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_373);
  gl_ram_g27658 : AO221D0BWP7T port map(A1 => gl_ram_n_120, A2 => gl_ram_n_84, B1 => gl_ram_n_200, B2 => FE_PHN219_gl_ram_ram_81_1, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_372);
  gl_ram_g27659 : AO221D0BWP7T port map(A1 => gl_ram_n_122, A2 => gl_ram_n_84, B1 => gl_ram_n_200, B2 => FE_PHN242_gl_ram_ram_81_2, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_371);
  gl_ram_g27660 : AO221D0BWP7T port map(A1 => gl_ram_n_114, A2 => gl_ram_n_108, B1 => gl_ram_n_227, B2 => FE_PHN605_gl_ram_ram_24_2, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_370);
  gl_ram_g27661 : AO221D0BWP7T port map(A1 => gl_ram_n_117, A2 => gl_ram_n_84, B1 => gl_ram_n_201, B2 => FE_PHN570_gl_ram_ram_82_0, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_369);
  gl_ram_g27662 : AO221D0BWP7T port map(A1 => gl_ram_n_116, A2 => gl_ram_n_84, B1 => gl_ram_n_201, B2 => FE_PHN408_gl_ram_ram_82_1, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_368);
  gl_ram_g27663 : AO221D0BWP7T port map(A1 => gl_ram_n_118, A2 => gl_ram_n_108, B1 => gl_ram_n_199, B2 => FE_PHN630_gl_ram_ram_25_0, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_367);
  gl_ram_g27664 : AO221D0BWP7T port map(A1 => gl_ram_n_85, A2 => gl_ram_n_84, B1 => gl_ram_n_201, B2 => FE_PHN294_gl_ram_ram_82_2, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_366);
  gl_ram_g27665 : AO221D0BWP7T port map(A1 => gl_ram_n_119, A2 => gl_ram_n_84, B1 => gl_ram_n_192, B2 => FE_PHN418_gl_ram_ram_83_0, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_365);
  gl_ram_g27666 : AO221D0BWP7T port map(A1 => gl_ram_n_120, A2 => gl_ram_n_108, B1 => gl_ram_n_199, B2 => FE_PHN423_gl_ram_ram_25_1, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_364);
  gl_ram_g27667 : AO221D0BWP7T port map(A1 => gl_ram_n_123, A2 => gl_ram_n_84, B1 => gl_ram_n_192, B2 => FE_PHN153_gl_ram_ram_83_1, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_363);
  gl_ram_g27668 : AO221D0BWP7T port map(A1 => gl_ram_n_121, A2 => gl_ram_n_84, B1 => gl_ram_n_192, B2 => FE_PHN188_gl_ram_ram_83_2, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_362);
  gl_ram_g27669 : AO221D0BWP7T port map(A1 => gl_ram_n_122, A2 => gl_ram_n_108, B1 => gl_ram_n_199, B2 => FE_PHN182_gl_ram_ram_25_2, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_361);
  gl_ram_g27670 : AO221D0BWP7T port map(A1 => gl_ram_n_133, A2 => gl_ram_n_84, B1 => gl_ram_n_222, B2 => FE_PHN154_gl_ram_ram_84_0, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_360);
  gl_ram_g27671 : AO221D0BWP7T port map(A1 => gl_ram_n_132, A2 => gl_ram_n_84, B1 => gl_ram_n_222, B2 => FE_PHN230_gl_ram_ram_84_1, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_359);
  gl_ram_g27672 : AO221D0BWP7T port map(A1 => gl_ram_n_117, A2 => gl_ram_n_108, B1 => gl_ram_n_197, B2 => FE_PHN176_gl_ram_ram_26_0, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_358);
  gl_ram_g27673 : AO221D0BWP7T port map(A1 => gl_ram_n_131, A2 => gl_ram_n_84, B1 => gl_ram_n_222, B2 => FE_PHN92_gl_ram_ram_84_2, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_357);
  gl_ram_g27674 : AO221D0BWP7T port map(A1 => gl_ram_n_86, A2 => gl_ram_n_113, B1 => gl_ram_n_217, B2 => FE_PHN553_gl_ram_ram_0_0, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_356);
  gl_ram_g27675 : AO221D0BWP7T port map(A1 => gl_ram_n_124, A2 => gl_ram_n_84, B1 => gl_ram_n_182, B2 => FE_PHN161_gl_ram_ram_85_0, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_355);
  gl_ram_g27676 : AO221D0BWP7T port map(A1 => gl_ram_n_116, A2 => gl_ram_n_108, B1 => gl_ram_n_197, B2 => FE_PHN223_gl_ram_ram_26_1, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_354);
  gl_ram_g27677 : AO221D0BWP7T port map(A1 => gl_ram_n_130, A2 => gl_ram_n_84, B1 => gl_ram_n_182, B2 => FE_PHN236_gl_ram_ram_85_1, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_353);
  gl_ram_g27678 : AO221D0BWP7T port map(A1 => gl_ram_n_87, A2 => gl_ram_n_84, B1 => gl_ram_n_182, B2 => FE_PHN109_gl_ram_ram_85_2, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_352);
  gl_ram_g27679 : AO221D0BWP7T port map(A1 => gl_ram_n_115, A2 => gl_ram_n_113, B1 => gl_ram_n_217, B2 => FE_PHN560_gl_ram_ram_0_1, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_351);
  gl_ram_g27680 : AO221D0BWP7T port map(A1 => gl_ram_n_134, A2 => gl_ram_n_84, B1 => gl_ram_n_152, B2 => FE_PHN291_gl_ram_ram_86_0, C => gl_ram_n_16, Z => gl_ram_n_350);
  gl_ram_g27681 : AO221D0BWP7T port map(A1 => gl_ram_n_85, A2 => gl_ram_n_108, B1 => gl_ram_n_197, B2 => FE_PHN218_gl_ram_ram_26_2, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_349);
  gl_ram_g27682 : AO221D0BWP7T port map(A1 => gl_ram_n_128, A2 => gl_ram_n_84, B1 => gl_ram_n_152, B2 => FE_PHN317_gl_ram_ram_86_1, C => gl_ram_n_16, Z => gl_ram_n_348);
  gl_ram_g27683 : AO221D0BWP7T port map(A1 => gl_ram_n_119, A2 => gl_ram_n_108, B1 => gl_ram_n_193, B2 => FE_PHN596_gl_ram_ram_27_0, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_347);
  gl_ram_g27684 : AO221D0BWP7T port map(A1 => gl_ram_n_127, A2 => gl_ram_n_84, B1 => gl_ram_n_152, B2 => FE_PHN298_gl_ram_ram_86_2, C => gl_ram_n_16, Z => gl_ram_n_346);
  gl_ram_g27685 : AO221D0BWP7T port map(A1 => gl_ram_n_126, A2 => gl_ram_n_84, B1 => gl_ram_n_184, B2 => FE_PHN112_gl_ram_ram_87_0, C => gl_ram_n_16, Z => gl_ram_n_345);
  gl_ram_g27686 : AO221D0BWP7T port map(A1 => gl_ram_n_123, A2 => gl_ram_n_108, B1 => gl_ram_n_193, B2 => FE_PHN555_gl_ram_ram_27_1, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_344);
  gl_ram_g27687 : AO221D0BWP7T port map(A1 => gl_ram_n_125, A2 => gl_ram_n_84, B1 => gl_ram_n_184, B2 => FE_PHN271_gl_ram_ram_87_1, C => gl_ram_n_16, Z => gl_ram_n_343);
  gl_ram_g27688 : AO221D0BWP7T port map(A1 => gl_ram_n_129, A2 => gl_ram_n_84, B1 => gl_ram_n_184, B2 => FE_PHN302_gl_ram_ram_87_2, C => gl_ram_n_16, Z => gl_ram_n_342);
  gl_ram_g27689 : AO221D0BWP7T port map(A1 => gl_ram_n_86, A2 => gl_ram_n_81, B1 => gl_ram_n_224, B2 => FE_PHN602_gl_ram_ram_88_0, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_341);
  gl_ram_g27690 : AO221D0BWP7T port map(A1 => gl_ram_n_121, A2 => gl_ram_n_108, B1 => gl_ram_n_193, B2 => FE_PHN635_gl_ram_ram_27_2, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_340);
  gl_ram_g27691 : AO221D0BWP7T port map(A1 => gl_ram_n_115, A2 => gl_ram_n_81, B1 => gl_ram_n_224, B2 => FE_PHN104_gl_ram_ram_88_1, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_339);
  gl_ram_g27692 : AO221D0BWP7T port map(A1 => gl_ram_n_133, A2 => gl_ram_n_108, B1 => gl_ram_n_220, B2 => FE_PHN251_gl_ram_ram_28_0, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_338);
  gl_ram_g27693 : AO221D0BWP7T port map(A1 => gl_ram_n_114, A2 => gl_ram_n_81, B1 => gl_ram_n_224, B2 => FE_PHN110_gl_ram_ram_88_2, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_337);
  gl_ram_g27694 : AO221D0BWP7T port map(A1 => gl_ram_n_118, A2 => gl_ram_n_81, B1 => gl_ram_n_196, B2 => FE_PHN624_gl_ram_ram_89_0, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_336);
  gl_ram_g27695 : AO221D0BWP7T port map(A1 => gl_ram_n_132, A2 => gl_ram_n_108, B1 => gl_ram_n_220, B2 => FE_PHN137_gl_ram_ram_28_1, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_335);
  gl_ram_g27696 : AO221D0BWP7T port map(A1 => gl_ram_n_120, A2 => gl_ram_n_81, B1 => gl_ram_n_196, B2 => FE_PHN216_gl_ram_ram_89_1, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_334);
  gl_ram_g27697 : AO221D0BWP7T port map(A1 => gl_ram_n_122, A2 => gl_ram_n_81, B1 => gl_ram_n_196, B2 => FE_PHN235_gl_ram_ram_89_2, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_333);
  gl_ram_g27698 : AO221D0BWP7T port map(A1 => gl_ram_n_131, A2 => gl_ram_n_108, B1 => gl_ram_n_220, B2 => FE_PHN151_gl_ram_ram_28_2, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_332);
  gl_ram_g27699 : AO221D0BWP7T port map(A1 => gl_ram_n_117, A2 => gl_ram_n_81, B1 => gl_ram_n_194, B2 => FE_PHN147_gl_ram_ram_90_0, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_331);
  gl_ram_g27700 : AO221D0BWP7T port map(A1 => gl_ram_n_114, A2 => gl_ram_n_113, B1 => gl_ram_n_217, B2 => FE_PHN523_gl_ram_ram_0_2, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_330);
  gl_ram_g27701 : AO221D0BWP7T port map(A1 => gl_ram_n_116, A2 => gl_ram_n_81, B1 => gl_ram_n_194, B2 => FE_PHN193_gl_ram_ram_90_1, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_329);
  gl_ram_g27702 : AO221D0BWP7T port map(A1 => gl_ram_n_124, A2 => gl_ram_n_108, B1 => gl_ram_n_148, B2 => FE_PHN119_gl_ram_ram_29_0, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_328);
  gl_ram_g27703 : AO221D0BWP7T port map(A1 => gl_ram_n_85, A2 => gl_ram_n_81, B1 => gl_ram_n_194, B2 => FE_PHN241_gl_ram_ram_90_2, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_327);
  gl_ram_g27704 : AO221D0BWP7T port map(A1 => gl_ram_n_119, A2 => gl_ram_n_81, B1 => gl_ram_n_190, B2 => FE_PHN168_gl_ram_ram_91_0, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_326);
  gl_ram_g27705 : AO221D0BWP7T port map(A1 => gl_ram_n_130, A2 => gl_ram_n_108, B1 => gl_ram_n_148, B2 => FE_PHN629_gl_ram_ram_29_1, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_325);
  gl_ram_g27706 : AO221D0BWP7T port map(A1 => gl_ram_n_123, A2 => gl_ram_n_81, B1 => gl_ram_n_190, B2 => FE_PHN574_gl_ram_ram_91_1, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_324);
  gl_ram_g27707 : AO221D0BWP7T port map(A1 => gl_ram_n_87, A2 => gl_ram_n_108, B1 => gl_ram_n_148, B2 => FE_PHN237_gl_ram_ram_29_2, C => FE_OFN38_gl_ram_n_16, Z => gl_ram_n_323);
  gl_ram_g27708 : AO221D0BWP7T port map(A1 => gl_ram_n_121, A2 => gl_ram_n_81, B1 => gl_ram_n_190, B2 => FE_PHN164_gl_ram_ram_91_2, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_322);
  gl_ram_g27709 : AO221D0BWP7T port map(A1 => gl_ram_n_118, A2 => gl_ram_n_113, B1 => gl_ram_n_163, B2 => FE_PHN561_gl_ram_ram_1_0, C => FE_OFN39_gl_ram_n_16, Z => gl_ram_n_321);
  gl_ram_g27710 : AO221D0BWP7T port map(A1 => gl_ram_n_133, A2 => gl_ram_n_81, B1 => gl_ram_n_219, B2 => FE_PHN159_gl_ram_ram_92_0, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_320);
  gl_ram_g27711 : AO221D0BWP7T port map(A1 => gl_ram_n_132, A2 => gl_ram_n_81, B1 => gl_ram_n_219, B2 => FE_PHN101_gl_ram_ram_92_1, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_319);
  gl_ram_g27712 : AO221D0BWP7T port map(A1 => gl_ram_n_134, A2 => gl_ram_n_108, B1 => gl_ram_n_153, B2 => FE_PHN201_gl_ram_ram_30_0, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_318);
  gl_ram_g27713 : AO221D0BWP7T port map(A1 => gl_ram_n_131, A2 => gl_ram_n_81, B1 => gl_ram_n_219, B2 => FE_PHN108_gl_ram_ram_92_2, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_317);
  gl_ram_g27714 : AO221D0BWP7T port map(A1 => gl_ram_n_124, A2 => gl_ram_n_81, B1 => gl_ram_n_185, B2 => FE_PHN220_gl_ram_ram_93_0, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_316);
  gl_ram_g27715 : AO221D0BWP7T port map(A1 => gl_ram_n_128, A2 => gl_ram_n_108, B1 => gl_ram_n_153, B2 => FE_PHN258_gl_ram_ram_30_1, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_315);
  gl_ram_g27716 : AO221D0BWP7T port map(A1 => gl_ram_n_130, A2 => gl_ram_n_81, B1 => gl_ram_n_185, B2 => FE_PHN190_gl_ram_ram_93_1, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_314);
  gl_ram_g27717 : AO222D0BWP7T port map(A1 => gl_ram_n_136, A2 => gl_ram_n_29, B1 => gl_ram_n_236, B2 => gl_ram_x_grid(2), C1 => gl_ram_n_188, C2 => gl_ram_n_2, Z => gl_ram_n_313);
  gl_ram_g27718 : AOI33D1BWP7T port map(A1 => gl_ram_n_230, A2 => gl_ram_n_47, A3 => gl_ram_y_grid(3), B1 => gl_ram_n_232, B2 => gl_ram_n_18, B3 => gl_ram_n_13, ZN => gl_ram_n_312);
  gl_ram_g27719 : MOAI22D0BWP7T port map(A1 => gl_ram_n_239, A2 => gl_ram_x_grid(3), B1 => gl_ram_n_235, B2 => gl_ram_n_21, ZN => gl_ram_n_311);
  gl_ram_g27720 : AO221D0BWP7T port map(A1 => gl_ram_n_115, A2 => gl_ram_n_50, B1 => gl_ram_n_103, B2 => FE_PHN114_gl_ram_ram_64_1, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_310);
  gl_ram_g27721 : AO221D0BWP7T port map(A1 => gl_ram_n_87, A2 => gl_ram_n_50, B1 => gl_ram_n_94, B2 => FE_PHN250_gl_ram_ram_69_2, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_309);
  gl_ram_g27722 : AO211D0BWP7T port map(A1 => gl_ram_ram_position(1), A2 => gl_ram_n_16, B => gl_ram_n_188, C => gl_ram_n_141, Z => gl_ram_n_308);
  gl_ram_g27723 : AO221D0BWP7T port map(A1 => gl_ram_n_86, A2 => gl_ram_n_51, B1 => gl_ram_n_107, B2 => FE_PHN210_gl_ram_ram_96_0, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_307);
  gl_ram_g27724 : AO221D0BWP7T port map(A1 => gl_ram_n_115, A2 => gl_ram_n_51, B1 => gl_ram_n_107, B2 => FE_PHN419_gl_ram_ram_96_1, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_306);
  gl_ram_g27725 : AO221D0BWP7T port map(A1 => gl_ram_n_114, A2 => gl_ram_n_51, B1 => gl_ram_n_107, B2 => FE_PHN426_gl_ram_ram_96_2, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_305);
  gl_ram_g27726 : AO221D0BWP7T port map(A1 => gl_ram_n_118, A2 => gl_ram_n_51, B1 => gl_ram_n_105, B2 => FE_PHN420_gl_ram_ram_97_0, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_304);
  gl_ram_g27727 : AO221D0BWP7T port map(A1 => gl_ram_n_120, A2 => gl_ram_n_51, B1 => gl_ram_n_105, B2 => FE_PHN650_gl_ram_ram_97_1, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_303);
  gl_ram_g27728 : AO221D0BWP7T port map(A1 => gl_ram_n_122, A2 => gl_ram_n_51, B1 => gl_ram_n_105, B2 => FE_PHN99_gl_ram_ram_97_2, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_302);
  gl_ram_g27729 : AO221D0BWP7T port map(A1 => gl_ram_n_117, A2 => gl_ram_n_51, B1 => gl_ram_n_104, B2 => FE_PHN257_gl_ram_ram_98_0, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_301);
  gl_ram_g27730 : AO221D0BWP7T port map(A1 => gl_ram_n_116, A2 => gl_ram_n_51, B1 => gl_ram_n_104, B2 => FE_PHN214_gl_ram_ram_98_1, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_300);
  gl_ram_g27731 : AO221D0BWP7T port map(A1 => gl_ram_n_85, A2 => gl_ram_n_51, B1 => gl_ram_n_104, B2 => FE_PHN409_gl_ram_ram_98_2, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_299);
  gl_ram_g27732 : AO221D0BWP7T port map(A1 => gl_ram_n_119, A2 => gl_ram_n_51, B1 => gl_ram_n_106, B2 => FE_PHN256_gl_ram_ram_99_0, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_298);
  gl_ram_g27733 : AO221D0BWP7T port map(A1 => gl_ram_n_123, A2 => gl_ram_n_51, B1 => gl_ram_n_106, B2 => FE_PHN248_gl_ram_ram_99_1, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_297);
  gl_ram_g27734 : AO221D0BWP7T port map(A1 => gl_ram_n_121, A2 => gl_ram_n_51, B1 => gl_ram_n_106, B2 => FE_PHN113_gl_ram_ram_99_2, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_296);
  gl_ram_g27735 : AO221D0BWP7T port map(A1 => gl_ram_n_86, A2 => gl_ram_n_50, B1 => gl_ram_n_103, B2 => FE_PHN221_gl_ram_ram_64_0, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_295);
  gl_ram_g27736 : AO221D0BWP7T port map(A1 => gl_ram_n_130, A2 => gl_ram_n_50, B1 => gl_ram_n_94, B2 => FE_PHN229_gl_ram_ram_69_1, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_294);
  gl_ram_g27737 : AO221D0BWP7T port map(A1 => gl_ram_n_114, A2 => gl_ram_n_50, B1 => gl_ram_n_103, B2 => FE_PHN252_gl_ram_ram_64_2, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_293);
  gl_ram_g27738 : AO221D0BWP7T port map(A1 => gl_ram_n_118, A2 => gl_ram_n_50, B1 => gl_ram_n_88, B2 => FE_PHN125_gl_ram_ram_65_0, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_292);
  gl_ram_g27739 : AO221D0BWP7T port map(A1 => gl_ram_n_120, A2 => gl_ram_n_50, B1 => gl_ram_n_88, B2 => FE_PHN144_gl_ram_ram_65_1, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_291);
  gl_ram_g27740 : AO221D0BWP7T port map(A1 => gl_ram_n_122, A2 => gl_ram_n_50, B1 => gl_ram_n_88, B2 => FE_PHN421_gl_ram_ram_65_2, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_290);
  gl_ram_g27741 : AO221D0BWP7T port map(A1 => gl_ram_n_117, A2 => gl_ram_n_50, B1 => gl_ram_n_89, B2 => FE_PHN416_gl_ram_ram_66_0, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_289);
  gl_ram_g27742 : AO221D0BWP7T port map(A1 => gl_ram_n_116, A2 => gl_ram_n_50, B1 => gl_ram_n_89, B2 => FE_PHN143_gl_ram_ram_66_1, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_288);
  gl_ram_g27743 : AO221D0BWP7T port map(A1 => gl_ram_n_85, A2 => gl_ram_n_50, B1 => gl_ram_n_89, B2 => FE_PHN280_gl_ram_ram_66_2, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_287);
  gl_ram_g27744 : AO221D0BWP7T port map(A1 => gl_ram_n_119, A2 => gl_ram_n_50, B1 => gl_ram_n_90, B2 => FE_PHN414_gl_ram_ram_67_0, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_286);
  gl_ram_g27745 : AO221D0BWP7T port map(A1 => gl_ram_n_123, A2 => gl_ram_n_50, B1 => gl_ram_n_90, B2 => FE_PHN200_gl_ram_ram_67_1, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_285);
  gl_ram_g27746 : AO221D0BWP7T port map(A1 => gl_ram_n_121, A2 => gl_ram_n_50, B1 => gl_ram_n_90, B2 => FE_PHN116_gl_ram_ram_67_2, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_284);
  gl_ram_g27747 : AO221D0BWP7T port map(A1 => gl_ram_n_133, A2 => gl_ram_n_50, B1 => gl_ram_n_97, B2 => FE_PHN264_gl_ram_ram_68_0, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_283);
  gl_ram_g27748 : AO221D0BWP7T port map(A1 => gl_ram_n_132, A2 => gl_ram_n_50, B1 => gl_ram_n_97, B2 => FE_PHN128_gl_ram_ram_68_1, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_282);
  gl_ram_g27749 : AO221D0BWP7T port map(A1 => gl_ram_n_131, A2 => gl_ram_n_50, B1 => gl_ram_n_97, B2 => FE_PHN103_gl_ram_ram_68_2, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_281);
  gl_ram_g27750 : AO221D0BWP7T port map(A1 => gl_ram_n_124, A2 => gl_ram_n_50, B1 => gl_ram_n_94, B2 => FE_PHN215_gl_ram_ram_69_0, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_280);
  gl_ram_g27753 : INVD0BWP7T port map(I => gl_ram_n_279, ZN => gl_ram_n_278);
  gl_ram_g27754 : AO221D0BWP7T port map(A1 => gl_ram_n_134, A2 => gl_ram_n_50, B1 => gl_ram_n_95, B2 => FE_PHN255_gl_ram_ram_70_0, C => gl_ram_n_16, Z => gl_ram_n_277);
  gl_ram_g27755 : AO221D0BWP7T port map(A1 => gl_ram_n_128, A2 => gl_ram_n_50, B1 => gl_ram_n_95, B2 => FE_PHN157_gl_ram_ram_70_1, C => gl_ram_n_16, Z => gl_ram_n_276);
  gl_ram_g27756 : AO221D0BWP7T port map(A1 => gl_ram_n_127, A2 => gl_ram_n_50, B1 => gl_ram_n_95, B2 => FE_PHN305_gl_ram_ram_70_2, C => gl_ram_n_16, Z => gl_ram_n_275);
  gl_ram_g27757 : AO221D0BWP7T port map(A1 => gl_ram_n_126, A2 => gl_ram_n_50, B1 => gl_ram_n_96, B2 => FE_PHN130_gl_ram_ram_71_0, C => gl_ram_n_16, Z => gl_ram_n_274);
  gl_ram_g27758 : AO221D0BWP7T port map(A1 => gl_ram_n_125, A2 => gl_ram_n_50, B1 => gl_ram_n_96, B2 => FE_PHN303_gl_ram_ram_71_1, C => gl_ram_n_16, Z => gl_ram_n_273);
  gl_ram_g27759 : AO221D0BWP7T port map(A1 => gl_ram_n_129, A2 => gl_ram_n_50, B1 => gl_ram_n_96, B2 => FE_PHN129_gl_ram_ram_71_2, C => gl_ram_n_16, Z => gl_ram_n_272);
  gl_ram_g27760 : AO221D0BWP7T port map(A1 => gl_ram_n_86, A2 => gl_ram_n_62, B1 => gl_ram_n_102, B2 => FE_PHN107_gl_ram_ram_72_0, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_271);
  gl_ram_g27761 : AO221D0BWP7T port map(A1 => gl_ram_n_115, A2 => gl_ram_n_62, B1 => gl_ram_n_102, B2 => FE_PHN139_gl_ram_ram_72_1, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_270);
  gl_ram_g27762 : AO221D0BWP7T port map(A1 => gl_ram_n_114, A2 => gl_ram_n_62, B1 => gl_ram_n_102, B2 => FE_PHN196_gl_ram_ram_72_2, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_269);
  gl_ram_g27763 : AO221D0BWP7T port map(A1 => gl_ram_n_118, A2 => gl_ram_n_62, B1 => gl_ram_n_91, B2 => FE_PHN417_gl_ram_ram_73_0, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_268);
  gl_ram_g27764 : AO221D0BWP7T port map(A1 => gl_ram_n_120, A2 => gl_ram_n_62, B1 => gl_ram_n_91, B2 => FE_PHN412_gl_ram_ram_73_1, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_267);
  gl_ram_g27765 : AO221D0BWP7T port map(A1 => gl_ram_n_122, A2 => gl_ram_n_62, B1 => gl_ram_n_91, B2 => FE_PHN604_gl_ram_ram_73_2, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_266);
  gl_ram_g27766 : AO221D0BWP7T port map(A1 => gl_ram_n_117, A2 => gl_ram_n_62, B1 => gl_ram_n_93, B2 => FE_PHN162_gl_ram_ram_74_0, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_265);
  gl_ram_g27767 : AO221D0BWP7T port map(A1 => gl_ram_n_116, A2 => gl_ram_n_62, B1 => gl_ram_n_93, B2 => FE_PHN246_gl_ram_ram_74_1, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_264);
  gl_ram_g27768 : AO221D0BWP7T port map(A1 => gl_ram_n_85, A2 => gl_ram_n_62, B1 => gl_ram_n_93, B2 => FE_PHN234_gl_ram_ram_74_2, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_263);
  gl_ram_g27769 : AO221D0BWP7T port map(A1 => gl_ram_n_119, A2 => gl_ram_n_62, B1 => gl_ram_n_92, B2 => FE_PHN580_gl_ram_ram_75_0, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_262);
  gl_ram_g27770 : AO221D0BWP7T port map(A1 => gl_ram_n_123, A2 => gl_ram_n_62, B1 => gl_ram_n_92, B2 => FE_PHN212_gl_ram_ram_75_1, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_261);
  gl_ram_g27771 : AO221D0BWP7T port map(A1 => gl_ram_n_121, A2 => gl_ram_n_62, B1 => gl_ram_n_92, B2 => FE_PHN191_gl_ram_ram_75_2, C => FE_OFN40_gl_ram_n_16, Z => gl_ram_n_260);
  gl_ram_g27772 : AO221D0BWP7T port map(A1 => gl_ram_n_133, A2 => gl_ram_n_62, B1 => gl_ram_n_98, B2 => FE_PHN286_gl_ram_ram_76_0, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_259);
  gl_ram_g27773 : AO221D0BWP7T port map(A1 => gl_ram_n_132, A2 => gl_ram_n_62, B1 => gl_ram_n_98, B2 => FE_PHN189_gl_ram_ram_76_1, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_258);
  gl_ram_g27774 : AO221D0BWP7T port map(A1 => gl_ram_n_131, A2 => gl_ram_n_62, B1 => gl_ram_n_98, B2 => FE_PHN270_gl_ram_ram_76_2, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_257);
  gl_ram_g27775 : AO221D0BWP7T port map(A1 => gl_ram_n_124, A2 => gl_ram_n_62, B1 => gl_ram_n_99, B2 => FE_PHN98_gl_ram_ram_77_0, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_256);
  gl_ram_g27776 : AO221D0BWP7T port map(A1 => gl_ram_n_130, A2 => gl_ram_n_62, B1 => gl_ram_n_99, B2 => FE_PHN199_gl_ram_ram_77_1, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_255);
  gl_ram_g27777 : AO221D0BWP7T port map(A1 => gl_ram_n_87, A2 => gl_ram_n_62, B1 => gl_ram_n_99, B2 => FE_PHN226_gl_ram_ram_77_2, C => FE_OFN37_gl_ram_n_16, Z => gl_ram_n_254);
  gl_ram_g27778 : AO221D0BWP7T port map(A1 => gl_ram_n_134, A2 => gl_ram_n_62, B1 => gl_ram_n_100, B2 => FE_PHN141_gl_ram_ram_78_0, C => gl_ram_n_16, Z => gl_ram_n_253);
  gl_ram_g27779 : AO221D0BWP7T port map(A1 => gl_ram_n_128, A2 => gl_ram_n_62, B1 => gl_ram_n_100, B2 => FE_PHN296_gl_ram_ram_78_1, C => gl_ram_n_16, Z => gl_ram_n_252);
  gl_ram_g27780 : AO221D0BWP7T port map(A1 => gl_ram_n_127, A2 => gl_ram_n_62, B1 => gl_ram_n_100, B2 => FE_PHN240_gl_ram_ram_78_2, C => gl_ram_n_16, Z => gl_ram_n_251);
  gl_ram_g27781 : AO221D0BWP7T port map(A1 => gl_ram_n_126, A2 => gl_ram_n_62, B1 => gl_ram_n_101, B2 => FE_PHN152_gl_ram_ram_79_0, C => gl_ram_n_16, Z => gl_ram_n_250);
  gl_ram_g27782 : AO221D0BWP7T port map(A1 => gl_ram_n_125, A2 => gl_ram_n_62, B1 => gl_ram_n_101, B2 => FE_PHN135_gl_ram_ram_79_1, C => gl_ram_n_16, Z => gl_ram_n_249);
  gl_ram_g27783 : AO221D0BWP7T port map(A1 => gl_ram_n_129, A2 => gl_ram_n_62, B1 => gl_ram_n_101, B2 => FE_PHN238_gl_ram_ram_79_2, C => gl_ram_n_16, Z => gl_ram_n_248);
  gl_ram_g27784 : OAI31D0BWP7T port map(A1 => sig_logic_y(2), A2 => gl_ram_n_9, A3 => gl_ram_n_69, B => gl_ram_n_238, ZN => gl_ram_n_247);
  gl_ram_g27785 : MAOI22D0BWP7T port map(A1 => gl_ram_n_230, A2 => gl_ram_y_grid(2), B1 => gl_ram_n_186, B2 => gl_ram_n_45, ZN => gl_ram_n_246);
  gl_ram_g27786 : AOI22D0BWP7T port map(A1 => gl_ram_n_136, A2 => gl_ram_n_28, B1 => gl_ram_n_233, B2 => gl_ram_x_grid(1), ZN => gl_ram_n_245);
  gl_ram_g27787 : OAI21D0BWP7T port map(A1 => gl_ram_n_135, A2 => gl_ram_n_8, B => gl_ram_n_242, ZN => gl_ram_n_279);
  gl_ram_g27788 : NR2D0BWP7T port map(A1 => gl_ram_n_234, A2 => gl_ram_x_grid(1), ZN => gl_ram_n_244);
  gl_ram_g27789 : IOA21D1BWP7T port map(A1 => gl_ram_n_76, A2 => sig_logic_y(0), B => gl_ram_n_143, ZN => gl_ram_n_243);
  gl_ram_g27793 : AOI22D0BWP7T port map(A1 => gl_ram_n_136, A2 => gl_ram_n_32, B1 => gl_ram_ram_position(2), B2 => gl_ram_n_16, ZN => gl_ram_n_241);
  gl_ram_g27794 : OAI222D0BWP7T port map(A1 => gl_ram_n_75, A2 => gl_ram_n_45, B1 => FE_PHN327_gl_ram_n_5, B2 => gl_ram_n_48, C1 => gl_ram_x_grid(3), C2 => gl_ram_n_21, ZN => gl_ram_n_240);
  gl_ram_g27795 : MAOI22D0BWP7T port map(A1 => gl_ram_n_136, A2 => gl_ram_n_14, B1 => gl_ram_n_137, B2 => gl_ram_y_grid(3), ZN => gl_ram_n_239);
  gl_ram_g27796 : AOI22D0BWP7T port map(A1 => gl_ram_n_139, A2 => gl_ram_n_9, B1 => gl_ram_y_grid(2), B2 => gl_ram_n_16, ZN => gl_ram_n_238);
  gl_ram_g27797 : OAI22D0BWP7T port map(A1 => gl_ram_n_138, A2 => gl_ram_n_9, B1 => gl_ram_n_4, B2 => gl_ram_n_15, ZN => gl_ram_n_237);
  gl_ram_g27798 : IND3D1BWP7T port map(A1 => gl_ram_n_135, B1 => gl_ram_x_grid(2), B2 => gl_ram_y_grid(0), ZN => gl_ram_n_242);
  gl_ram_g27799 : CKND1BWP7T port map(I => gl_ram_n_233, ZN => gl_ram_n_234);
  gl_ram_g27800 : INVD1BWP7T port map(I => gl_ram_n_231, ZN => gl_ram_n_232);
  gl_ram_g27802 : NR2D0BWP7T port map(A1 => gl_ram_n_135, A2 => gl_ram_y_grid(0), ZN => gl_ram_n_236);
  gl_ram_g27803 : AN2D0BWP7T port map(A1 => gl_ram_n_136, A2 => gl_ram_n_4, Z => gl_ram_n_235);
  gl_ram_g27804 : NR2D1BWP7T port map(A1 => gl_ram_n_135, A2 => gl_ram_x_grid(2), ZN => gl_ram_n_233);
  gl_ram_g27805 : ND2D1BWP7T port map(A1 => gl_ram_n_136, A2 => gl_ram_y_grid(3), ZN => gl_ram_n_231);
  gl_ram_g27806 : NR2D1BWP7T port map(A1 => gl_ram_n_135, A2 => gl_ram_n_12, ZN => gl_ram_n_230);
  gl_ram_g27807 : ND2D1BWP7T port map(A1 => gl_ram_n_56, A2 => gl_ram_n_109, ZN => gl_ram_n_229);
  gl_ram_g27808 : ND2D1BWP7T port map(A1 => gl_ram_n_57, A2 => gl_ram_n_109, ZN => gl_ram_n_228);
  gl_ram_g27809 : ND2D1BWP7T port map(A1 => gl_ram_n_55, A2 => gl_ram_n_108, ZN => gl_ram_n_227);
  gl_ram_g27810 : ND2D1BWP7T port map(A1 => gl_ram_n_55, A2 => gl_ram_n_112, ZN => gl_ram_n_226);
  gl_ram_g27811 : ND2D1BWP7T port map(A1 => gl_ram_n_55, A2 => gl_ram_n_84, ZN => gl_ram_n_225);
  gl_ram_g27812 : ND2D1BWP7T port map(A1 => gl_ram_n_55, A2 => gl_ram_n_81, ZN => gl_ram_n_224);
  gl_ram_g27813 : ND2D1BWP7T port map(A1 => gl_ram_n_55, A2 => gl_ram_n_83, ZN => gl_ram_n_223);
  gl_ram_g27814 : ND2D1BWP7T port map(A1 => gl_ram_n_59, A2 => gl_ram_n_84, ZN => gl_ram_n_222);
  gl_ram_g27815 : ND2D1BWP7T port map(A1 => gl_ram_n_59, A2 => gl_ram_n_112, ZN => gl_ram_n_221);
  gl_ram_g27816 : ND2D1BWP7T port map(A1 => gl_ram_n_59, A2 => gl_ram_n_108, ZN => gl_ram_n_220);
  gl_ram_g27817 : ND2D1BWP7T port map(A1 => gl_ram_n_59, A2 => gl_ram_n_81, ZN => gl_ram_n_219);
  gl_ram_g27818 : ND2D1BWP7T port map(A1 => gl_ram_n_55, A2 => gl_ram_n_111, ZN => gl_ram_n_218);
  gl_ram_g27819 : ND2D1BWP7T port map(A1 => gl_ram_n_55, A2 => gl_ram_n_113, ZN => gl_ram_n_217);
  gl_ram_g27820 : ND2D1BWP7T port map(A1 => gl_ram_n_59, A2 => gl_ram_n_83, ZN => gl_ram_n_216);
  gl_ram_g27821 : ND2D1BWP7T port map(A1 => gl_ram_n_55, A2 => gl_ram_n_110, ZN => gl_ram_n_215);
  gl_ram_g27822 : ND2D1BWP7T port map(A1 => gl_ram_n_55, A2 => gl_ram_n_82, ZN => gl_ram_n_214);
  gl_ram_g27823 : ND2D1BWP7T port map(A1 => gl_ram_n_55, A2 => gl_ram_n_109, ZN => gl_ram_n_213);
  gl_ram_g27824 : ND2D1BWP7T port map(A1 => gl_ram_n_58, A2 => gl_ram_n_110, ZN => gl_ram_n_212);
  gl_ram_g27825 : ND2D1BWP7T port map(A1 => gl_ram_n_56, A2 => gl_ram_n_110, ZN => gl_ram_n_211);
  gl_ram_g27826 : ND2D1BWP7T port map(A1 => gl_ram_n_57, A2 => gl_ram_n_110, ZN => gl_ram_n_210);
  gl_ram_g27827 : ND2D1BWP7T port map(A1 => gl_ram_n_58, A2 => gl_ram_n_82, ZN => gl_ram_n_209);
  gl_ram_g27828 : ND2D1BWP7T port map(A1 => gl_ram_n_57, A2 => gl_ram_n_82, ZN => gl_ram_n_208);
  gl_ram_g27829 : ND2D1BWP7T port map(A1 => gl_ram_n_56, A2 => gl_ram_n_82, ZN => gl_ram_n_207);
  gl_ram_g27830 : ND2D1BWP7T port map(A1 => gl_ram_n_59, A2 => gl_ram_n_111, ZN => gl_ram_n_206);
  gl_ram_g27831 : ND2D1BWP7T port map(A1 => gl_ram_n_59, A2 => gl_ram_n_113, ZN => gl_ram_n_205);
  gl_ram_g27832 : ND2D1BWP7T port map(A1 => gl_ram_n_59, A2 => gl_ram_n_82, ZN => gl_ram_n_204);
  gl_ram_g27833 : ND2D1BWP7T port map(A1 => gl_ram_n_59, A2 => gl_ram_n_110, ZN => gl_ram_n_203);
  gl_ram_g27834 : ND2D1BWP7T port map(A1 => gl_ram_n_59, A2 => gl_ram_n_109, ZN => gl_ram_n_202);
  gl_ram_g27835 : ND2D1BWP7T port map(A1 => gl_ram_n_52, A2 => gl_ram_n_84, ZN => gl_ram_n_201);
  gl_ram_g27836 : ND2D1BWP7T port map(A1 => gl_ram_n_54, A2 => gl_ram_n_84, ZN => gl_ram_n_200);
  gl_ram_g27837 : ND2D1BWP7T port map(A1 => gl_ram_n_54, A2 => gl_ram_n_108, ZN => gl_ram_n_199);
  gl_ram_g27838 : ND2D1BWP7T port map(A1 => gl_ram_n_54, A2 => gl_ram_n_112, ZN => gl_ram_n_198);
  gl_ram_g27839 : ND2D1BWP7T port map(A1 => gl_ram_n_52, A2 => gl_ram_n_108, ZN => gl_ram_n_197);
  gl_ram_g27840 : ND2D1BWP7T port map(A1 => gl_ram_n_54, A2 => gl_ram_n_81, ZN => gl_ram_n_196);
  gl_ram_g27841 : ND2D1BWP7T port map(A1 => gl_ram_n_52, A2 => gl_ram_n_112, ZN => gl_ram_n_195);
  gl_ram_g27842 : ND2D1BWP7T port map(A1 => gl_ram_n_52, A2 => gl_ram_n_81, ZN => gl_ram_n_194);
  gl_ram_g27843 : ND2D1BWP7T port map(A1 => gl_ram_n_53, A2 => gl_ram_n_108, ZN => gl_ram_n_193);
  gl_ram_g27844 : ND2D1BWP7T port map(A1 => gl_ram_n_53, A2 => gl_ram_n_84, ZN => gl_ram_n_192);
  gl_ram_g27845 : ND2D1BWP7T port map(A1 => gl_ram_n_53, A2 => gl_ram_n_112, ZN => gl_ram_n_191);
  gl_ram_g27846 : ND2D1BWP7T port map(A1 => gl_ram_n_53, A2 => gl_ram_n_81, ZN => gl_ram_n_190);
  gl_ram_g27847 : ND2D1BWP7T port map(A1 => gl_ram_n_58, A2 => gl_ram_n_109, ZN => gl_ram_n_189);
  gl_ram_g27850 : OAI22D0BWP7T port map(A1 => gl_ram_n_60, A2 => FE_PHN464_sig_logic_y_0, B1 => FE_PHN327_gl_ram_n_5, B2 => gl_ram_n_15, ZN => gl_ram_n_146);
  gl_ram_g27851 : OAI22D0BWP7T port map(A1 => gl_ram_n_49, A2 => gl_ram_n_41, B1 => gl_ram_n_2, B2 => gl_ram_n_15, ZN => gl_ram_n_145);
  gl_ram_g27852 : OAI22D0BWP7T port map(A1 => gl_ram_n_21, A2 => gl_ram_n_45, B1 => gl_ram_n_46, B2 => gl_ram_y_grid(0), ZN => gl_ram_n_144);
  gl_ram_g27853 : AOI22D0BWP7T port map(A1 => gl_ram_n_70, A2 => gl_ram_n_9, B1 => gl_ram_y_grid(1), B2 => gl_ram_n_16, ZN => gl_ram_n_143);
  gl_ram_g27854 : AO22D0BWP7T port map(A1 => gl_ram_n_61, A2 => gl_ram_x_grid(0), B1 => gl_ram_n_16, B2 => gl_ram_ram_position(0), Z => gl_ram_n_142);
  gl_ram_g27855 : NR3D0BWP7T port map(A1 => gl_ram_n_60, A2 => gl_ram_y_grid(0), A3 => gl_ram_n_3, ZN => gl_ram_n_141);
  gl_ram_g27856 : IND3D1BWP7T port map(A1 => gl_ram_n_135, B1 => gl_ram_n_12, B2 => gl_ram_n_45, ZN => gl_ram_n_140);
  gl_ram_g27857 : NR3D0BWP7T port map(A1 => gl_ram_n_60, A2 => FE_PHN327_gl_ram_n_5, A3 => gl_ram_x_grid(1), ZN => gl_ram_n_188);
  gl_ram_g27858 : NR3D0BWP7T port map(A1 => gl_ram_n_60, A2 => gl_ram_n_4, A3 => gl_ram_y_grid(2), ZN => gl_ram_n_187);
  gl_ram_g27859 : OA21D0BWP7T port map(A1 => gl_ram_n_60, A2 => gl_ram_n_21, B => gl_ram_n_135, Z => gl_ram_n_186);
  gl_ram_g27860 : ND2D1BWP7T port map(A1 => gl_ram_n_57, A2 => gl_ram_n_81, ZN => gl_ram_n_185);
  gl_ram_g27861 : ND2D1BWP7T port map(A1 => gl_ram_n_58, A2 => gl_ram_n_84, ZN => gl_ram_n_184);
  gl_ram_g27862 : ND2D1BWP7T port map(A1 => gl_ram_n_58, A2 => gl_ram_n_112, ZN => gl_ram_n_183);
  gl_ram_g27863 : ND2D1BWP7T port map(A1 => gl_ram_n_57, A2 => gl_ram_n_84, ZN => gl_ram_n_182);
  gl_ram_g27864 : ND2D1BWP7T port map(A1 => gl_ram_n_54, A2 => gl_ram_n_83, ZN => gl_ram_n_181);
  gl_ram_g27865 : ND2D1BWP7T port map(A1 => gl_ram_n_52, A2 => gl_ram_n_83, ZN => gl_ram_n_180);
  gl_ram_g27866 : ND2D1BWP7T port map(A1 => gl_ram_n_53, A2 => gl_ram_n_83, ZN => gl_ram_n_179);
  gl_ram_g27867 : ND2D1BWP7T port map(A1 => gl_ram_n_58, A2 => gl_ram_n_113, ZN => gl_ram_n_178);
  gl_ram_g27868 : ND2D1BWP7T port map(A1 => gl_ram_n_58, A2 => gl_ram_n_111, ZN => gl_ram_n_177);
  gl_ram_g27869 : ND2D1BWP7T port map(A1 => gl_ram_n_58, A2 => gl_ram_n_83, ZN => gl_ram_n_176);
  gl_ram_g27870 : ND2D1BWP7T port map(A1 => gl_ram_n_57, A2 => gl_ram_n_113, ZN => gl_ram_n_175);
  gl_ram_g27871 : ND2D1BWP7T port map(A1 => gl_ram_n_56, A2 => gl_ram_n_113, ZN => gl_ram_n_174);
  gl_ram_g27872 : ND2D1BWP7T port map(A1 => gl_ram_n_57, A2 => gl_ram_n_83, ZN => gl_ram_n_173);
  gl_ram_g27873 : ND2D1BWP7T port map(A1 => gl_ram_n_56, A2 => gl_ram_n_83, ZN => gl_ram_n_172);
  gl_ram_g27874 : ND2D1BWP7T port map(A1 => gl_ram_n_57, A2 => gl_ram_n_111, ZN => gl_ram_n_171);
  gl_ram_g27875 : ND2D1BWP7T port map(A1 => gl_ram_n_56, A2 => gl_ram_n_111, ZN => gl_ram_n_170);
  gl_ram_g27876 : ND2D1BWP7T port map(A1 => gl_ram_n_54, A2 => gl_ram_n_82, ZN => gl_ram_n_169);
  gl_ram_g27877 : ND2D1BWP7T port map(A1 => gl_ram_n_52, A2 => gl_ram_n_82, ZN => gl_ram_n_168);
  gl_ram_g27878 : ND2D1BWP7T port map(A1 => gl_ram_n_53, A2 => gl_ram_n_82, ZN => gl_ram_n_167);
  gl_ram_g27879 : ND2D1BWP7T port map(A1 => gl_ram_n_52, A2 => gl_ram_n_113, ZN => gl_ram_n_166);
  gl_ram_g27880 : ND2D1BWP7T port map(A1 => gl_ram_n_52, A2 => gl_ram_n_111, ZN => gl_ram_n_165);
  gl_ram_g27881 : ND2D1BWP7T port map(A1 => gl_ram_n_54, A2 => gl_ram_n_111, ZN => gl_ram_n_164);
  gl_ram_g27882 : ND2D1BWP7T port map(A1 => gl_ram_n_54, A2 => gl_ram_n_113, ZN => gl_ram_n_163);
  gl_ram_g27883 : ND2D1BWP7T port map(A1 => gl_ram_n_53, A2 => gl_ram_n_113, ZN => gl_ram_n_162);
  gl_ram_g27884 : ND2D1BWP7T port map(A1 => gl_ram_n_53, A2 => gl_ram_n_111, ZN => gl_ram_n_161);
  gl_ram_g27885 : ND2D1BWP7T port map(A1 => gl_ram_n_53, A2 => gl_ram_n_109, ZN => gl_ram_n_160);
  gl_ram_g27886 : ND2D1BWP7T port map(A1 => gl_ram_n_52, A2 => gl_ram_n_109, ZN => gl_ram_n_159);
  gl_ram_g27887 : ND2D1BWP7T port map(A1 => gl_ram_n_54, A2 => gl_ram_n_109, ZN => gl_ram_n_158);
  gl_ram_g27888 : ND2D1BWP7T port map(A1 => gl_ram_n_54, A2 => gl_ram_n_110, ZN => gl_ram_n_157);
  gl_ram_g27889 : ND2D1BWP7T port map(A1 => gl_ram_n_58, A2 => gl_ram_n_81, ZN => gl_ram_n_156);
  gl_ram_g27890 : ND2D1BWP7T port map(A1 => gl_ram_n_57, A2 => gl_ram_n_112, ZN => gl_ram_n_155);
  gl_ram_g27891 : ND2D1BWP7T port map(A1 => gl_ram_n_56, A2 => gl_ram_n_81, ZN => gl_ram_n_154);
  gl_ram_g27892 : ND2D1BWP7T port map(A1 => gl_ram_n_56, A2 => gl_ram_n_108, ZN => gl_ram_n_153);
  gl_ram_g27893 : ND2D1BWP7T port map(A1 => gl_ram_n_56, A2 => gl_ram_n_84, ZN => gl_ram_n_152);
  gl_ram_g27894 : ND2D1BWP7T port map(A1 => gl_ram_n_56, A2 => gl_ram_n_112, ZN => gl_ram_n_151);
  gl_ram_g27895 : ND2D1BWP7T port map(A1 => gl_ram_n_53, A2 => gl_ram_n_110, ZN => gl_ram_n_150);
  gl_ram_g27896 : ND2D1BWP7T port map(A1 => gl_ram_n_52, A2 => gl_ram_n_110, ZN => gl_ram_n_149);
  gl_ram_g27897 : ND2D1BWP7T port map(A1 => gl_ram_n_57, A2 => gl_ram_n_108, ZN => gl_ram_n_148);
  gl_ram_g27898 : ND2D1BWP7T port map(A1 => gl_ram_n_58, A2 => gl_ram_n_108, ZN => gl_ram_n_147);
  gl_ram_g27899 : INVD0BWP7T port map(I => gl_ram_n_138, ZN => gl_ram_n_139);
  gl_ram_g27900 : ND2D1BWP7T port map(A1 => gl_ram_n_70, A2 => sig_logic_y(2), ZN => gl_ram_n_138);
  gl_ram_g27901 : ND2D1BWP7T port map(A1 => gl_ram_n_61, A2 => gl_ram_n_12, ZN => gl_ram_n_137);
  gl_ram_g27902 : NR2D1BWP7T port map(A1 => gl_ram_n_60, A2 => gl_ram_y_grid(1), ZN => gl_ram_n_136);
  gl_ram_g27903 : ND2D1BWP7T port map(A1 => gl_ram_n_61, A2 => gl_ram_y_grid(1), ZN => gl_ram_n_135);
  gl_ram_g27904 : NR2XD0BWP7T port map(A1 => gl_ram_n_65, A2 => gl_ram_n_36, ZN => gl_ram_n_134);
  gl_ram_g27905 : NR2XD0BWP7T port map(A1 => gl_ram_n_65, A2 => gl_ram_n_33, ZN => gl_ram_n_133);
  gl_ram_g27906 : NR2XD0BWP7T port map(A1 => gl_ram_n_66, A2 => gl_ram_n_33, ZN => gl_ram_n_132);
  gl_ram_g27907 : NR2XD0BWP7T port map(A1 => gl_ram_n_64, A2 => gl_ram_n_33, ZN => gl_ram_n_131);
  gl_ram_g27908 : NR2XD0BWP7T port map(A1 => gl_ram_n_66, A2 => gl_ram_n_35, ZN => gl_ram_n_130);
  gl_ram_g27909 : NR2XD0BWP7T port map(A1 => gl_ram_n_64, A2 => gl_ram_n_34, ZN => gl_ram_n_129);
  gl_ram_g27910 : NR2XD0BWP7T port map(A1 => gl_ram_n_66, A2 => gl_ram_n_36, ZN => gl_ram_n_128);
  gl_ram_g27911 : NR2XD0BWP7T port map(A1 => gl_ram_n_64, A2 => gl_ram_n_36, ZN => gl_ram_n_127);
  gl_ram_g27912 : NR2XD0BWP7T port map(A1 => gl_ram_n_65, A2 => gl_ram_n_34, ZN => gl_ram_n_126);
  gl_ram_g27913 : NR2XD0BWP7T port map(A1 => gl_ram_n_66, A2 => gl_ram_n_34, ZN => gl_ram_n_125);
  gl_ram_g27914 : NR2XD0BWP7T port map(A1 => gl_ram_n_65, A2 => gl_ram_n_35, ZN => gl_ram_n_124);
  gl_ram_g27915 : NR2XD0BWP7T port map(A1 => gl_ram_n_67, A2 => gl_ram_n_34, ZN => gl_ram_n_123);
  gl_ram_g27916 : NR2XD0BWP7T port map(A1 => gl_ram_n_68, A2 => gl_ram_n_35, ZN => gl_ram_n_122);
  gl_ram_g27917 : NR2XD0BWP7T port map(A1 => gl_ram_n_68, A2 => gl_ram_n_34, ZN => gl_ram_n_121);
  gl_ram_g27918 : NR2XD0BWP7T port map(A1 => gl_ram_n_67, A2 => gl_ram_n_35, ZN => gl_ram_n_120);
  gl_ram_g27919 : NR2XD0BWP7T port map(A1 => gl_ram_n_63, A2 => gl_ram_n_34, ZN => gl_ram_n_119);
  gl_ram_g27920 : NR2XD0BWP7T port map(A1 => gl_ram_n_63, A2 => gl_ram_n_35, ZN => gl_ram_n_118);
  gl_ram_g27921 : NR2XD0BWP7T port map(A1 => gl_ram_n_63, A2 => gl_ram_n_36, ZN => gl_ram_n_117);
  gl_ram_g27922 : NR2XD0BWP7T port map(A1 => gl_ram_n_67, A2 => gl_ram_n_36, ZN => gl_ram_n_116);
  gl_ram_g27923 : NR2XD0BWP7T port map(A1 => gl_ram_n_67, A2 => gl_ram_n_33, ZN => gl_ram_n_115);
  gl_ram_g27924 : NR2XD0BWP7T port map(A1 => gl_ram_n_68, A2 => gl_ram_n_33, ZN => gl_ram_n_114);
  gl_ram_g27925 : CKAN2D1BWP7T port map(A1 => gl_ram_n_74, A2 => gl_ram_n_0, Z => gl_ram_n_113);
  gl_ram_g27926 : CKAN2D1BWP7T port map(A1 => gl_ram_n_74, A2 => gl_ram_ram_position(4), Z => gl_ram_n_112);
  gl_ram_g27927 : CKAN2D1BWP7T port map(A1 => gl_ram_n_71, A2 => gl_ram_n_0, Z => gl_ram_n_111);
  gl_ram_g27928 : NR2D1P5BWP7T port map(A1 => gl_ram_n_72, A2 => gl_ram_ram_position(4), ZN => gl_ram_n_110);
  gl_ram_g27929 : NR2D1P5BWP7T port map(A1 => gl_ram_n_72, A2 => gl_ram_n_0, ZN => gl_ram_n_109);
  gl_ram_g27930 : CKAN2D1BWP7T port map(A1 => gl_ram_n_71, A2 => gl_ram_ram_position(4), Z => gl_ram_n_108);
  gl_ram_g27931 : OAI22D0BWP7T port map(A1 => gl_ram_n_38, A2 => gl_ram_n_41, B1 => gl_ram_n_1, B2 => gl_ram_n_15, ZN => FE_PHN365_gl_ram_n_80);
  gl_ram_g27932 : OAI22D0BWP7T port map(A1 => gl_ram_n_45, A2 => gl_ram_y_grid(3), B1 => gl_ram_n_4, B2 => gl_ram_x_grid(3), ZN => gl_ram_n_79);
  gl_ram_g27933 : OAI22D0BWP7T port map(A1 => gl_ram_n_31, A2 => gl_ram_n_41, B1 => gl_ram_n_3, B2 => gl_ram_n_15, ZN => gl_ram_n_78);
  gl_ram_g27934 : OAI31D0BWP7T port map(A1 => sig_logic_x(0), A2 => gl_ram_n_25, A3 => gl_ram_n_41, B => gl_ram_n_20, ZN => gl_ram_n_77);
  gl_ram_g27935 : OA211D0BWP7T port map(A1 => sig_logic_y(3), A2 => sig_logic_y(2), B => gl_ram_n_37, C => sig_logic_y(1), Z => gl_ram_n_76);
  gl_ram_g27936 : ND2D1BWP7T port map(A1 => gl_ram_n_55, A2 => gl_ram_n_51, ZN => gl_ram_n_107);
  gl_ram_g27937 : ND2D1BWP7T port map(A1 => gl_ram_n_53, A2 => gl_ram_n_51, ZN => gl_ram_n_106);
  gl_ram_g27938 : ND2D1BWP7T port map(A1 => gl_ram_n_54, A2 => gl_ram_n_51, ZN => gl_ram_n_105);
  gl_ram_g27939 : ND2D1BWP7T port map(A1 => gl_ram_n_52, A2 => gl_ram_n_51, ZN => gl_ram_n_104);
  gl_ram_g27940 : ND2D1BWP7T port map(A1 => gl_ram_n_55, A2 => gl_ram_n_50, ZN => gl_ram_n_103);
  gl_ram_g27941 : ND2D1BWP7T port map(A1 => gl_ram_n_55, A2 => gl_ram_n_62, ZN => gl_ram_n_102);
  gl_ram_g27942 : ND2D1BWP7T port map(A1 => gl_ram_n_58, A2 => gl_ram_n_62, ZN => gl_ram_n_101);
  gl_ram_g27943 : ND2D1BWP7T port map(A1 => gl_ram_n_56, A2 => gl_ram_n_62, ZN => gl_ram_n_100);
  gl_ram_g27944 : ND2D1BWP7T port map(A1 => gl_ram_n_57, A2 => gl_ram_n_62, ZN => gl_ram_n_99);
  gl_ram_g27945 : ND2D1BWP7T port map(A1 => gl_ram_n_59, A2 => gl_ram_n_62, ZN => gl_ram_n_98);
  gl_ram_g27946 : ND2D1BWP7T port map(A1 => gl_ram_n_59, A2 => gl_ram_n_50, ZN => gl_ram_n_97);
  gl_ram_g27947 : ND2D1BWP7T port map(A1 => gl_ram_n_58, A2 => gl_ram_n_50, ZN => gl_ram_n_96);
  gl_ram_g27948 : ND2D1BWP7T port map(A1 => gl_ram_n_56, A2 => gl_ram_n_50, ZN => gl_ram_n_95);
  gl_ram_g27949 : ND2D1BWP7T port map(A1 => gl_ram_n_57, A2 => gl_ram_n_50, ZN => gl_ram_n_94);
  gl_ram_g27950 : ND2D1BWP7T port map(A1 => gl_ram_n_52, A2 => gl_ram_n_62, ZN => gl_ram_n_93);
  gl_ram_g27951 : ND2D1BWP7T port map(A1 => gl_ram_n_53, A2 => gl_ram_n_62, ZN => gl_ram_n_92);
  gl_ram_g27952 : ND2D1BWP7T port map(A1 => gl_ram_n_54, A2 => gl_ram_n_62, ZN => gl_ram_n_91);
  gl_ram_g27953 : ND2D1BWP7T port map(A1 => gl_ram_n_53, A2 => gl_ram_n_50, ZN => gl_ram_n_90);
  gl_ram_g27954 : ND2D1BWP7T port map(A1 => gl_ram_n_52, A2 => gl_ram_n_50, ZN => gl_ram_n_89);
  gl_ram_g27955 : ND2D1BWP7T port map(A1 => gl_ram_n_54, A2 => gl_ram_n_50, ZN => gl_ram_n_88);
  gl_ram_g27956 : NR2XD0BWP7T port map(A1 => gl_ram_n_64, A2 => gl_ram_n_35, ZN => gl_ram_n_87);
  gl_ram_g27957 : NR2XD0BWP7T port map(A1 => gl_ram_n_63, A2 => gl_ram_n_33, ZN => gl_ram_n_86);
  gl_ram_g27958 : NR2XD0BWP7T port map(A1 => gl_ram_n_68, A2 => gl_ram_n_36, ZN => gl_ram_n_85);
  gl_ram_g27959 : AN3D1BWP7T port map(A1 => gl_ram_n_42, A2 => gl_ram_ram_position(4), A3 => gl_ram_ram_position(6), Z => gl_ram_n_84);
  gl_ram_g27960 : NR2D1P5BWP7T port map(A1 => gl_ram_n_73, A2 => gl_ram_n_0, ZN => gl_ram_n_83);
  gl_ram_g27961 : NR2D1P5BWP7T port map(A1 => gl_ram_n_73, A2 => gl_ram_ram_position(4), ZN => gl_ram_n_82);
  gl_ram_g27962 : AN3D1BWP7T port map(A1 => gl_ram_n_43, A2 => gl_ram_ram_position(4), A3 => gl_ram_ram_position(6), Z => gl_ram_n_81);
  gl_ram_g27963 : INVD0BWP7T port map(I => gl_ram_n_21, ZN => gl_ram_n_75);
  gl_ram_g27964 : INVD1BWP7T port map(I => gl_ram_n_69, ZN => gl_ram_n_70);
  gl_ram_g27965 : INR2XD0BWP7T port map(A1 => gl_ram_n_42, B1 => gl_ram_ram_position(6), ZN => gl_ram_n_74);
  gl_ram_g27966 : IND2D1BWP7T port map(A1 => gl_ram_ram_position(3), B1 => gl_ram_n_44, ZN => gl_ram_n_73);
  gl_ram_g27967 : ND2D1BWP7T port map(A1 => gl_ram_n_44, A2 => gl_ram_ram_position(3), ZN => gl_ram_n_72);
  gl_ram_g27968 : INR2XD0BWP7T port map(A1 => gl_ram_n_43, B1 => gl_ram_ram_position(6), ZN => gl_ram_n_71);
  gl_ram_g27969 : ND2D1BWP7T port map(A1 => gl_ram_n_37, A2 => sig_logic_y(3), ZN => gl_ram_n_69);
  gl_ram_g27970 : ND2D1BWP7T port map(A1 => sig_output_color(2), A2 => gl_ram_n_40, ZN => gl_ram_n_68);
  gl_ram_g27971 : ND2D1BWP7T port map(A1 => gl_ram_n_40, A2 => sig_output_color(1), ZN => gl_ram_n_67);
  gl_ram_g27972 : ND2D1BWP7T port map(A1 => gl_ram_n_39, A2 => sig_output_color(1), ZN => gl_ram_n_66);
  gl_ram_g27973 : ND2D1BWP7T port map(A1 => gl_ram_n_39, A2 => sig_output_color(0), ZN => gl_ram_n_65);
  gl_ram_g27974 : ND2D1BWP7T port map(A1 => sig_output_color(2), A2 => gl_ram_n_39, ZN => gl_ram_n_64);
  gl_ram_g27975 : ND2D1BWP7T port map(A1 => gl_ram_n_40, A2 => sig_output_color(0), ZN => gl_ram_n_63);
  gl_ram_g27976 : INR2D2BWP7T port map(A1 => gl_ram_n_43, B1 => gl_ram_n_10, ZN => gl_ram_n_62);
  gl_ram_g27977 : INVD1BWP7T port map(I => gl_ram_n_61, ZN => gl_ram_n_60);
  gl_ram_g27978 : AOI22D0BWP7T port map(A1 => gl_ram_n_24, A2 => sig_logic_x(3), B1 => gl_ram_n_17, B2 => sig_logic_x(2), ZN => gl_ram_n_49);
  gl_ram_g27979 : NR2D1BWP7T port map(A1 => gl_ram_n_41, A2 => gl_ram_n_27, ZN => gl_ram_n_61);
  gl_ram_g27980 : INR2XD0BWP7T port map(A1 => gl_ram_n_39, B1 => gl_ram_n_33, ZN => gl_ram_n_59);
  gl_ram_g27981 : INR2XD0BWP7T port map(A1 => gl_ram_n_39, B1 => gl_ram_n_34, ZN => gl_ram_n_58);
  gl_ram_g27982 : INR2XD0BWP7T port map(A1 => gl_ram_n_39, B1 => gl_ram_n_35, ZN => gl_ram_n_57);
  gl_ram_g27983 : INR2XD0BWP7T port map(A1 => gl_ram_n_39, B1 => gl_ram_n_36, ZN => gl_ram_n_56);
  gl_ram_g27984 : INR2XD0BWP7T port map(A1 => gl_ram_n_40, B1 => gl_ram_n_33, ZN => gl_ram_n_55);
  gl_ram_g27985 : INR2XD0BWP7T port map(A1 => gl_ram_n_40, B1 => gl_ram_n_35, ZN => gl_ram_n_54);
  gl_ram_g27986 : INR2XD0BWP7T port map(A1 => gl_ram_n_40, B1 => gl_ram_n_34, ZN => gl_ram_n_53);
  gl_ram_g27987 : INR2XD0BWP7T port map(A1 => gl_ram_n_40, B1 => gl_ram_n_36, ZN => gl_ram_n_52);
  gl_ram_g27988 : NR3D1BWP7T port map(A1 => gl_ram_n_10, A2 => gl_ram_n_23, A3 => gl_ram_ram_position(3), ZN => gl_ram_n_51);
  gl_ram_g27989 : INR2D2BWP7T port map(A1 => gl_ram_n_42, B1 => gl_ram_n_10, ZN => gl_ram_n_50);
  gl_ram_g27990 : INVD0BWP7T port map(I => gl_ram_n_47, ZN => gl_ram_n_48);
  gl_ram_g27991 : INVD1BWP7T port map(I => gl_ram_n_46, ZN => gl_ram_n_45);
  gl_ram_g27992 : HA1D0BWP7T port map(A => gl_ram_x_grid(3), B => gl_ram_y_grid(2), CO => gl_ram_n_46, S => gl_ram_n_47);
  gl_ram_g27993 : IND2D1BWP7T port map(A1 => gl_ram_n_24, B1 => sig_logic_x(3), ZN => gl_ram_n_38);
  gl_ram_g27994 : NR2XD0BWP7T port map(A1 => gl_ram_n_23, A2 => gl_ram_ram_position(6), ZN => gl_ram_n_44);
  gl_ram_g27995 : CKAN2D1BWP7T port map(A1 => gl_ram_n_30, A2 => gl_ram_ram_position(3), Z => gl_ram_n_43);
  gl_ram_g27996 : INR2XD0BWP7T port map(A1 => gl_ram_n_30, B1 => gl_ram_ram_position(3), ZN => gl_ram_n_42);
  gl_ram_g27997 : OR2D1BWP7T port map(A1 => gl_ram_n_22, A2 => gl_ram_n_16, Z => gl_ram_n_41);
  gl_ram_g27998 : NR2XD0BWP7T port map(A1 => gl_ram_n_22, A2 => gl_ram_ram_position(2), ZN => gl_ram_n_40);
  gl_ram_g27999 : INR2XD0BWP7T port map(A1 => gl_ram_ram_position(2), B1 => gl_ram_n_22, ZN => gl_ram_n_39);
  gl_ram_g28000 : OAI22D0BWP7T port map(A1 => gl_ram_n_8, A2 => gl_ram_x_grid(2), B1 => gl_ram_n_7, B2 => gl_ram_n_2, ZN => gl_ram_n_32);
  gl_ram_g28001 : MAOI22D0BWP7T port map(A1 => sig_logic_x(0), A2 => sig_logic_x(1), B1 => gl_ram_n_17, B2 => gl_ram_n_11, ZN => gl_ram_n_31);
  gl_ram_g28002 : NR2XD0BWP7T port map(A1 => gl_ram_n_27, A2 => gl_ram_n_16, ZN => gl_ram_n_37);
  gl_ram_g28003 : IND3D1BWP7T port map(A1 => gl_ram_ram_position(0), B1 => gl_ram_ram_position(1), B2 => gl_ram_n_26, ZN => gl_ram_n_36);
  gl_ram_g28004 : IND3D1BWP7T port map(A1 => gl_ram_ram_position(1), B1 => gl_ram_ram_position(0), B2 => gl_ram_n_26, ZN => gl_ram_n_35);
  gl_ram_g28005 : ND3D0BWP7T port map(A1 => gl_ram_n_26, A2 => gl_ram_ram_position(0), A3 => gl_ram_ram_position(1), ZN => gl_ram_n_34);
  gl_ram_g28006 : OR3D1BWP7T port map(A1 => gl_ram_ram_position(0), A2 => gl_ram_ram_position(1), A3 => gl_ram_n_27, Z => gl_ram_n_33);
  gl_ram_g28007 : INVD0BWP7T port map(I => gl_ram_n_28, ZN => gl_ram_n_29);
  gl_ram_g28008 : INVD1BWP7T port map(I => gl_ram_n_27, ZN => gl_ram_n_26);
  gl_ram_g28009 : INR2D1BWP7T port map(A1 => gl_ram_n_11, B1 => sig_logic_x(1), ZN => gl_ram_n_25);
  gl_ram_g28010 : NR2XD0BWP7T port map(A1 => gl_ram_ram_position(5), A2 => gl_ram_n_19, ZN => gl_ram_n_30);
  gl_ram_g28011 : ND2D1BWP7T port map(A1 => gl_ram_n_13, A2 => gl_ram_y_grid(0), ZN => gl_ram_n_28);
  gl_ram_g28012 : INR2XD0BWP7T port map(A1 => gl_ram_n_11, B1 => gl_ram_n_17, ZN => gl_ram_n_27);
  gl_ram_g28013 : ND2D1BWP7T port map(A1 => gl_ram_x_grid(0), A2 => gl_ram_n_16, ZN => gl_ram_n_20);
  gl_ram_g28014 : NR2XD0BWP7T port map(A1 => gl_ram_n_17, A2 => sig_logic_x(2), ZN => gl_ram_n_24);
  gl_ram_g28015 : IND2D1BWP7T port map(A1 => gl_ram_n_19, B1 => gl_ram_ram_position(5), ZN => gl_ram_n_23);
  gl_ram_g28016 : AOI21D0BWP7T port map(A1 => sig_logic_y(1), A2 => sig_logic_y(2), B => sig_logic_y(3), ZN => gl_ram_n_22);
  gl_ram_g28017 : ND2D1BWP7T port map(A1 => gl_ram_n_7, A2 => gl_ram_x_grid(2), ZN => gl_ram_n_21);
  gl_ram_g28018 : INVD1BWP7T port map(I => gl_ram_n_16, ZN => gl_ram_n_15);
  gl_ram_g28019 : ND2D0BWP7T port map(A1 => gl_ram_y_grid(0), A2 => gl_ram_y_grid(3), ZN => gl_ram_n_14);
  gl_ram_g28020 : ND2D1BWP7T port map(A1 => sig_rescount, A2 => sig_draw, ZN => gl_ram_n_19);
  gl_ram_g28021 : NR2D0BWP7T port map(A1 => gl_ram_y_grid(2), A2 => gl_ram_x_grid(3), ZN => gl_ram_n_18);
  gl_ram_g28022 : OR2D1BWP7T port map(A1 => sig_logic_x(0), A2 => sig_logic_x(1), Z => gl_ram_n_17);
  gl_ram_g28023 : OR2D2BWP7T port map(A1 => FE_OFN35_reset, A2 => sig_middelsteknop, Z => gl_ram_n_16);
  gl_ram_g28024 : INVD0BWP7T port map(I => gl_ram_n_8, ZN => gl_ram_n_7);
  gl_ram_g28025 : ND2D1BWP7T port map(A1 => gl_ram_x_grid(2), A2 => gl_ram_x_grid(1), ZN => gl_ram_n_13);
  gl_ram_g28026 : NR2XD0BWP7T port map(A1 => gl_ram_x_grid(2), A2 => gl_ram_y_grid(0), ZN => gl_ram_n_12);
  gl_ram_g28027 : NR2XD0BWP7T port map(A1 => sig_logic_x(2), A2 => sig_logic_x(3), ZN => gl_ram_n_11);
  gl_ram_g28028 : ND2D1BWP7T port map(A1 => gl_ram_n_0, A2 => gl_ram_ram_position(6), ZN => gl_ram_n_10);
  gl_ram_g28029 : NR2XD0BWP7T port map(A1 => sig_logic_y(0), A2 => sig_logic_y(1), ZN => gl_ram_n_9);
  gl_ram_g28030 : CKND2D1BWP7T port map(A1 => gl_ram_x_grid(1), A2 => gl_ram_y_grid(0), ZN => gl_ram_n_8);
  gl_ram_ram_position_reg_4 : DFD1BWP7T port map(CP => CTS_23, D => FE_PHN366_gl_ram_n_568, Q => gl_ram_ram_position(4), QN => gl_ram_n_0);
  gl_ram_x_grid_reg_1 : DFD1BWP7T port map(CP => CTS_19, D => FE_PHN361_gl_ram_n_78, Q => gl_ram_x_grid(1), QN => gl_ram_n_3);
  gl_ram_x_grid_reg_2 : DFD1BWP7T port map(CP => CTS_19, D => FE_PHN392_gl_ram_n_145, Q => gl_ram_x_grid(2), QN => gl_ram_n_2);
  gl_ram_x_grid_reg_3 : DFD1BWP7T port map(CP => CTS_19, D => gl_ram_n_80, Q => gl_ram_x_grid(3), QN => gl_ram_n_1);
  gl_ram_y_grid_reg_0 : DFD1BWP7T port map(CP => CTS_19, D => gl_ram_n_146, Q => gl_ram_y_grid(0), QN => gl_ram_n_5);
  gl_ram_y_grid_reg_2 : DFD1BWP7T port map(CP => CTS_19, D => FE_PHN377_gl_ram_n_247, Q => gl_ram_y_grid(2), QN => gl_ram_n_6);
  gl_ram_y_grid_reg_3 : DFD1BWP7T port map(CP => CTS_19, D => FE_PHN369_gl_ram_n_237, Q => gl_ram_y_grid(3), QN => gl_ram_n_4);
  gl_gr_lg_lcountdown_g204 : NR3D0BWP7T port map(A1 => gl_gr_lg_lcountdown_n_29, A2 => gl_gr_lg_lcountdown_n_22, A3 => gl_gr_lg_lcountdown_n_23, ZN => sig_countlow);
  gl_gr_lg_lcountdown_g205 : ND3D0BWP7T port map(A1 => gl_gr_lg_sig_countdown(10), A2 => gl_gr_lg_sig_countdown(9), A3 => FE_PHN353_gl_gr_lg_sig_countdown_0, ZN => gl_gr_lg_lcountdown_n_23);
  gl_gr_lg_lcountdown_g206 : ND4D0BWP7T port map(A1 => FE_PHN354_gl_gr_lg_sig_countdown_2, A2 => FE_PHN352_gl_gr_lg_sig_countdown_1, A3 => FE_PHN319_gl_gr_lg_sig_countdown_3, A4 => gl_gr_lg_sig_countdown(8), ZN => gl_gr_lg_lcountdown_n_22);
  gl_gr_lg_lcountdown_g207 : ND4D0BWP7T port map(A1 => FE_PHN355_gl_gr_lg_sig_countdown_5, A2 => gl_gr_lg_sig_countdown(4), A3 => gl_gr_lg_sig_countdown(6), A4 => gl_gr_lg_sig_countdown(7), ZN => gl_gr_lg_lcountdown_n_29);
  gl_gr_lg_lcountdown_count_c_reg_7 : DFKCNQD1BWP7T port map(CN => gl_gr_lg_lcountdown_n_1, CP => CTS_19, D => FE_PHN399_gl_gr_lg_lcountdown_n_21, Q => gl_gr_lg_sig_countdown(7));
  gl_gr_lg_lcountdown_count_c_reg_10 : DFKCNQD1BWP7T port map(CN => gl_gr_lg_lcountdown_n_1, CP => CTS_19, D => FE_PHN401_gl_gr_lg_lcountdown_n_20, Q => FE_PHN356_gl_gr_lg_sig_countdown_10);
  gl_gr_lg_lcountdown_g458 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_lcountdown_n_18, A2 => gl_gr_lg_sig_countdown(7), B1 => gl_gr_lg_lcountdown_n_18, B2 => gl_gr_lg_sig_countdown(7), ZN => gl_gr_lg_lcountdown_n_21);
  gl_gr_lg_lcountdown_count_c_reg_6 : DFKCNQD1BWP7T port map(CN => gl_gr_lg_lcountdown_n_1, CP => CTS_19, D => FE_PHN403_gl_gr_lg_lcountdown_n_19, Q => gl_gr_lg_sig_countdown(6));
  gl_gr_lg_lcountdown_count_c_reg_9 : DFKCNQD1BWP7T port map(CN => gl_gr_lg_lcountdown_n_1, CP => CTS_19, D => FE_PHN404_gl_gr_lg_lcountdown_n_17, Q => gl_gr_lg_sig_countdown(9));
  gl_gr_lg_lcountdown_g461 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_lcountdown_n_16, A2 => gl_gr_lg_sig_countdown(10), B1 => gl_gr_lg_lcountdown_n_16, B2 => gl_gr_lg_sig_countdown(10), ZN => gl_gr_lg_lcountdown_n_20);
  gl_gr_lg_lcountdown_count_c_reg_5 : DFKCNQD1BWP7T port map(CN => gl_gr_lg_lcountdown_n_1, CP => CTS_19, D => FE_PHN435_gl_gr_lg_lcountdown_n_15, Q => gl_gr_lg_sig_countdown(5));
  gl_gr_lg_lcountdown_g463 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_lcountdown_n_14, A2 => gl_gr_lg_sig_countdown(6), B1 => gl_gr_lg_lcountdown_n_14, B2 => gl_gr_lg_sig_countdown(6), ZN => gl_gr_lg_lcountdown_n_19);
  gl_gr_lg_lcountdown_g464 : IND2D1BWP7T port map(A1 => gl_gr_lg_lcountdown_n_14, B1 => gl_gr_lg_sig_countdown(6), ZN => gl_gr_lg_lcountdown_n_18);
  gl_gr_lg_lcountdown_count_c_reg_8 : DFKCNQD1BWP7T port map(CN => gl_gr_lg_lcountdown_n_1, CP => CTS_19, D => FE_PHN405_gl_gr_lg_lcountdown_n_13, Q => gl_gr_lg_sig_countdown(8));
  gl_gr_lg_lcountdown_g466 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_lcountdown_n_12, A2 => gl_gr_lg_sig_countdown(9), B1 => gl_gr_lg_lcountdown_n_12, B2 => gl_gr_lg_sig_countdown(9), ZN => gl_gr_lg_lcountdown_n_17);
  gl_gr_lg_lcountdown_count_c_reg_4 : DFKCNQD1BWP7T port map(CN => gl_gr_lg_lcountdown_n_1, CP => CTS_19, D => gl_gr_lg_lcountdown_n_11, Q => gl_gr_lg_sig_countdown(4));
  gl_gr_lg_lcountdown_g468 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_lcountdown_n_9, A2 => FE_PHN355_gl_gr_lg_sig_countdown_5, B1 => gl_gr_lg_lcountdown_n_9, B2 => FE_PHN355_gl_gr_lg_sig_countdown_5, ZN => gl_gr_lg_lcountdown_n_15);
  gl_gr_lg_lcountdown_g469 : IND2D1BWP7T port map(A1 => gl_gr_lg_lcountdown_n_12, B1 => gl_gr_lg_sig_countdown(9), ZN => gl_gr_lg_lcountdown_n_16);
  gl_gr_lg_lcountdown_g470 : IND2D1BWP7T port map(A1 => gl_gr_lg_lcountdown_n_9, B1 => FE_PHN355_gl_gr_lg_sig_countdown_5, ZN => gl_gr_lg_lcountdown_n_14);
  gl_gr_lg_lcountdown_g471 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_lcountdown_n_10, A2 => gl_gr_lg_sig_countdown(8), B1 => gl_gr_lg_lcountdown_n_10, B2 => gl_gr_lg_sig_countdown(8), ZN => gl_gr_lg_lcountdown_n_13);
  gl_gr_lg_lcountdown_count_c_reg_3 : DFKCNQD1BWP7T port map(CN => gl_gr_lg_lcountdown_n_1, CP => CTS_19, D => FE_PHN402_gl_gr_lg_lcountdown_n_8, Q => gl_gr_lg_sig_countdown(3));
  gl_gr_lg_lcountdown_g473 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_lcountdown_n_7, A2 => gl_gr_lg_sig_countdown(4), B1 => gl_gr_lg_lcountdown_n_7, B2 => gl_gr_lg_sig_countdown(4), ZN => FE_PHN400_gl_gr_lg_lcountdown_n_11);
  gl_gr_lg_lcountdown_g474 : IND2D1BWP7T port map(A1 => gl_gr_lg_lcountdown_n_10, B1 => gl_gr_lg_sig_countdown(8), ZN => gl_gr_lg_lcountdown_n_12);
  gl_gr_lg_lcountdown_g475 : OR2D1BWP7T port map(A1 => gl_gr_lg_lcountdown_n_7, A2 => gl_gr_lg_lcountdown_n_29, Z => gl_gr_lg_lcountdown_n_10);
  gl_gr_lg_lcountdown_g476 : IND2D1BWP7T port map(A1 => gl_gr_lg_lcountdown_n_7, B1 => gl_gr_lg_sig_countdown(4), ZN => gl_gr_lg_lcountdown_n_9);
  gl_gr_lg_lcountdown_count_c_reg_2 : DFKCNQD1BWP7T port map(CN => gl_gr_lg_lcountdown_n_1, CP => CTS_19, D => gl_gr_lg_lcountdown_n_6, Q => gl_gr_lg_sig_countdown(2));
  gl_gr_lg_lcountdown_g478 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_lcountdown_n_5, A2 => FE_PHN319_gl_gr_lg_sig_countdown_3, B1 => gl_gr_lg_lcountdown_n_5, B2 => FE_PHN319_gl_gr_lg_sig_countdown_3, ZN => gl_gr_lg_lcountdown_n_8);
  gl_gr_lg_lcountdown_g479 : IND2D1BWP7T port map(A1 => gl_gr_lg_lcountdown_n_5, B1 => FE_PHN319_gl_gr_lg_sig_countdown_3, ZN => gl_gr_lg_lcountdown_n_7);
  gl_gr_lg_lcountdown_count_c_reg_1 : DFKCNQD1BWP7T port map(CN => gl_gr_lg_lcountdown_n_1, CP => CTS_19, D => FE_PHN443_gl_gr_lg_lcountdown_n_4, Q => gl_gr_lg_sig_countdown(1));
  gl_gr_lg_lcountdown_g481 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_lcountdown_n_3, A2 => FE_PHN354_gl_gr_lg_sig_countdown_2, B1 => gl_gr_lg_lcountdown_n_3, B2 => FE_PHN354_gl_gr_lg_sig_countdown_2, ZN => gl_gr_lg_lcountdown_n_6);
  gl_gr_lg_lcountdown_g482 : IND2D1BWP7T port map(A1 => gl_gr_lg_lcountdown_n_3, B1 => FE_PHN354_gl_gr_lg_sig_countdown_2, ZN => gl_gr_lg_lcountdown_n_5);
  gl_gr_lg_lcountdown_count_c_reg_0 : DFKCNQD1BWP7T port map(CN => gl_gr_lg_lcountdown_n_1, CP => CTS_19, D => gl_gr_lg_lcountdown_n_2, Q => gl_gr_lg_sig_countdown(0));
  gl_gr_lg_lcountdown_g484 : MOAI22D0BWP7T port map(A1 => FE_PHN398_gl_gr_lg_lcountdown_n_0, A2 => FE_PHN352_gl_gr_lg_sig_countdown_1, B1 => FE_PHN398_gl_gr_lg_lcountdown_n_0, B2 => FE_PHN352_gl_gr_lg_sig_countdown_1, ZN => gl_gr_lg_lcountdown_n_4);
  gl_gr_lg_lcountdown_g485 : IND2D1BWP7T port map(A1 => FE_PHN398_gl_gr_lg_lcountdown_n_0, B1 => FE_PHN352_gl_gr_lg_sig_countdown_1, ZN => gl_gr_lg_lcountdown_n_3);
  gl_gr_lg_lcountdown_g486 : CKXOR2D1BWP7T port map(A1 => FE_PHN353_gl_gr_lg_sig_countdown_0, A2 => FE_PHN396_gl_gr_lg_lcountdown_sig_edge_fall, Z => FE_PHN445_gl_gr_lg_lcountdown_n_2);
  gl_gr_lg_lcountdown_g487 : NR2D1BWP7T port map(A1 => FE_OFN35_reset, A2 => sig_middelsteknop, ZN => gl_gr_lg_lcountdown_n_1);
  gl_gr_lg_lcountdown_g488 : ND2D1BWP7T port map(A1 => FE_PHN353_gl_gr_lg_sig_countdown_0, A2 => FE_PHN396_gl_gr_lg_lcountdown_sig_edge_fall, ZN => gl_gr_lg_lcountdown_n_0);
  gl_gr_lg_lcountdown_l_edge_g12 : NR2XD0BWP7T port map(A1 => gl_gr_lg_lcountdown_l_edge_reg2, A2 => FE_PHN304_gl_gr_lg_lcountdown_l_edge_reg1, ZN => gl_gr_lg_lcountdown_sig_edge_fall);
  gl_gr_lg_lcountdown_l_edge_reg2_reg : DFD0BWP7T port map(CP => CTS_19, D => FE_PHN304_gl_gr_lg_lcountdown_l_edge_reg1, Q => UNCONNECTED, QN => gl_gr_lg_lcountdown_l_edge_reg2);
  gl_gr_lg_lcountdown_l_edge_reg1_reg : DFQD1BWP7T port map(CP => CTS_19, D => FE_PHN362_gl_sig_v, Q => gl_gr_lg_lcountdown_l_edge_reg1);
  gl_vga_buf_G1_Q_reg : EDFQD1BWP7T port map(CP => CTS_20, D => gl_Gint, E => FE_DBTN0_reset, Q => gl_vga_buf_Gint);
  gl_vga_buf_G2_Q_reg : EDFQD0BWP7T port map(CP => CTS_20, D => FE_PHN67_gl_vga_buf_Gint, E => FE_DBTN0_reset, Q => FE_OFN32_G);
  gl_vga_buf_V1_Q_reg : EDFQD0BWP7T port map(CP => CTS_19, D => FE_PHN362_gl_sig_v, E => FE_DBTN0_reset, Q => FE_PHN88_gl_vga_buf_Vint);
  gl_vga_buf_V2_Q_reg : EDFQD0BWP7T port map(CP => CTS_19, D => gl_vga_buf_Vint, E => FE_DBTN0_reset, Q => FE_OFN30_V);
  gl_vga_buf_H1_Q_reg : EDFQD0BWP7T port map(CP => CTS_19, D => gl_Hint, E => FE_DBTN0_reset, Q => gl_vga_buf_Hint);
  gl_vga_buf_H2_Q_reg : EDFQD0BWP7T port map(CP => CTS_20, D => FE_PHN70_gl_vga_buf_Hint, E => FE_DBTN0_reset, Q => FE_OFN31_H);
  gl_vga_buf_B1_Q_reg : EDFQD1BWP7T port map(CP => CTS_20, D => gl_Bint, E => FE_DBTN0_reset, Q => gl_vga_buf_Bint);
  gl_gr_lg_le_g56 : INVD0BWP7T port map(I => gl_gr_lg_le_n_32, ZN => gl_gr_lg_le_n_31);
  gl_gr_lg_le_g447 : AN4D1BWP7T port map(A1 => gl_gr_lg_le_n_29, A2 => gl_gr_lg_le_n_28, A3 => gl_gr_lg_le_n_26, A4 => gl_gr_lg_le_n_21, Z => gl_gr_lg_le_n_32);
  gl_gr_lg_le_g448 : NR4D0BWP7T port map(A1 => gl_gr_lg_le_n_22, A2 => gl_gr_lg_le_n_27, A3 => gl_gr_lg_le_n_25, A4 => gl_gr_lg_le_n_20, ZN => gl_gr_lg_le_n_29);
  gl_gr_lg_le_g449 : NR2XD0BWP7T port map(A1 => gl_gr_lg_le_n_24, A2 => gl_gr_lg_le_n_23, ZN => gl_gr_lg_le_n_28);
  gl_gr_lg_le_g450 : CKXOR2D0BWP7T port map(A1 => sig_logic_x(1), A2 => gl_gr_lg_local_x(1), Z => gl_gr_lg_le_n_27);
  gl_gr_lg_le_g451 : MOAI22D0BWP7T port map(A1 => sig_logic_y(3), A2 => gl_gr_lg_local_y(3), B1 => sig_logic_y(3), B2 => gl_gr_lg_local_y(3), ZN => gl_gr_lg_le_n_26);
  gl_gr_lg_le_g452 : CKXOR2D0BWP7T port map(A1 => sig_logic_x(2), A2 => gl_gr_lg_local_x(2), Z => gl_gr_lg_le_n_25);
  gl_gr_lg_le_g453 : MAOI22D0BWP7T port map(A1 => sig_logic_y(2), A2 => gl_gr_lg_local_y(2), B1 => sig_logic_y(2), B2 => gl_gr_lg_local_y(2), ZN => gl_gr_lg_le_n_24);
  gl_gr_lg_le_g454 : MAOI22D0BWP7T port map(A1 => sig_logic_y(1), A2 => gl_gr_lg_local_y(1), B1 => sig_logic_y(1), B2 => gl_gr_lg_local_y(1), ZN => gl_gr_lg_le_n_23);
  gl_gr_lg_le_g455 : CKXOR2D0BWP7T port map(A1 => sig_logic_x(0), A2 => gl_gr_lg_local_x(0), Z => gl_gr_lg_le_n_22);
  gl_gr_lg_le_g456 : MOAI22D0BWP7T port map(A1 => sig_logic_y(0), A2 => gl_gr_lg_local_y(0), B1 => sig_logic_y(0), B2 => gl_gr_lg_local_y(0), ZN => gl_gr_lg_le_n_21);
  gl_gr_lg_le_g457 : CKXOR2D0BWP7T port map(A1 => sig_logic_x(3), A2 => gl_gr_lg_local_x(3), Z => gl_gr_lg_le_n_20);
  gl_gr_lg_le_new_count_e_reg_9 : LNQD1BWP7T port map(D => gl_gr_lg_le_n_19, EN => gl_gr_lg_le_n_18, Q => gl_gr_lg_le_new_count_e(9));
  gl_gr_lg_le_g342 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_le_n_16, A2 => gl_sig_e(9), B1 => gl_gr_lg_le_n_16, B2 => gl_sig_e(9), ZN => gl_gr_lg_le_n_19);
  gl_gr_lg_le_new_count_e_reg_8 : LNQD1BWP7T port map(D => gl_gr_lg_le_n_17, EN => gl_gr_lg_le_n_18, Q => gl_gr_lg_le_new_count_e(8));
  gl_gr_lg_le_g344 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_le_n_14, A2 => gl_sig_e(8), B1 => gl_gr_lg_le_n_14, B2 => gl_sig_e(8), ZN => gl_gr_lg_le_n_17);
  gl_gr_lg_le_new_count_e_reg_7 : LNQD1BWP7T port map(D => gl_gr_lg_le_n_15, EN => gl_gr_lg_le_n_18, Q => gl_gr_lg_le_new_count_e(7));
  gl_gr_lg_le_g346 : IND2D1BWP7T port map(A1 => gl_gr_lg_le_n_14, B1 => gl_sig_e(8), ZN => gl_gr_lg_le_n_16);
  gl_gr_lg_le_g347 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_le_n_12, A2 => gl_sig_e(7), B1 => gl_gr_lg_le_n_12, B2 => gl_sig_e(7), ZN => gl_gr_lg_le_n_15);
  gl_gr_lg_le_new_count_e_reg_6 : LNQD1BWP7T port map(D => gl_gr_lg_le_n_13, EN => gl_gr_lg_le_n_18, Q => gl_gr_lg_le_new_count_e(6));
  gl_gr_lg_le_g349 : IND2D1BWP7T port map(A1 => gl_gr_lg_le_n_12, B1 => gl_sig_e(7), ZN => gl_gr_lg_le_n_14);
  gl_gr_lg_le_g350 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_le_n_10, A2 => gl_sig_e(6), B1 => gl_gr_lg_le_n_10, B2 => gl_sig_e(6), ZN => gl_gr_lg_le_n_13);
  gl_gr_lg_le_new_count_e_reg_5 : LNQD1BWP7T port map(D => gl_gr_lg_le_n_11, EN => gl_gr_lg_le_n_18, Q => gl_gr_lg_le_new_count_e(5));
  gl_gr_lg_le_g352 : IND2D1BWP7T port map(A1 => gl_gr_lg_le_n_10, B1 => gl_sig_e(6), ZN => gl_gr_lg_le_n_12);
  gl_gr_lg_le_g353 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_le_n_8, A2 => gl_sig_e(5), B1 => gl_gr_lg_le_n_8, B2 => gl_sig_e(5), ZN => gl_gr_lg_le_n_11);
  gl_gr_lg_le_new_count_e_reg_4 : LNQD1BWP7T port map(D => gl_gr_lg_le_n_9, EN => gl_gr_lg_le_n_18, Q => gl_gr_lg_le_new_count_e(4));
  gl_gr_lg_le_g355 : IND2D1BWP7T port map(A1 => gl_gr_lg_le_n_8, B1 => gl_sig_e(5), ZN => gl_gr_lg_le_n_10);
  gl_gr_lg_le_g356 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_le_n_6, A2 => gl_sig_e(4), B1 => gl_gr_lg_le_n_6, B2 => gl_sig_e(4), ZN => gl_gr_lg_le_n_9);
  gl_gr_lg_le_new_count_e_reg_3 : LNQD1BWP7T port map(D => gl_gr_lg_le_n_7, EN => gl_gr_lg_le_n_18, Q => gl_gr_lg_le_new_count_e(3));
  gl_gr_lg_le_g358 : IND2D1BWP7T port map(A1 => gl_gr_lg_le_n_6, B1 => gl_sig_e(4), ZN => gl_gr_lg_le_n_8);
  gl_gr_lg_le_g359 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_le_n_4, A2 => gl_sig_e(3), B1 => gl_gr_lg_le_n_4, B2 => gl_sig_e(3), ZN => gl_gr_lg_le_n_7);
  gl_gr_lg_le_new_count_e_reg_2 : LNQD1BWP7T port map(D => gl_gr_lg_le_n_5, EN => gl_gr_lg_le_n_18, Q => gl_gr_lg_le_new_count_e(2));
  gl_gr_lg_le_g361 : IND2D1BWP7T port map(A1 => gl_gr_lg_le_n_4, B1 => gl_sig_e(3), ZN => gl_gr_lg_le_n_6);
  gl_gr_lg_le_g362 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_le_n_2, A2 => gl_sig_e(2), B1 => gl_gr_lg_le_n_2, B2 => gl_sig_e(2), ZN => gl_gr_lg_le_n_5);
  gl_gr_lg_le_new_count_e_reg_1 : LNQD1BWP7T port map(D => gl_gr_lg_le_n_3, EN => gl_gr_lg_le_n_18, Q => FE_PHN49_gl_gr_lg_le_new_count_e_1);
  gl_gr_lg_le_g364 : IND2D1BWP7T port map(A1 => gl_gr_lg_le_n_2, B1 => gl_sig_e(2), ZN => gl_gr_lg_le_n_4);
  gl_gr_lg_le_g365 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_le_n_0, A2 => gl_sig_e(1), B1 => gl_gr_lg_le_n_0, B2 => gl_sig_e(1), ZN => gl_gr_lg_le_n_3);
  gl_gr_lg_le_new_count_e_reg_0 : LNQD1BWP7T port map(D => gl_gr_lg_le_n_1, EN => gl_gr_lg_le_n_18, Q => FE_PHN50_gl_gr_lg_le_new_count_e_0);
  gl_gr_lg_le_g367 : IND2D1BWP7T port map(A1 => gl_gr_lg_le_n_0, B1 => gl_sig_e(1), ZN => gl_gr_lg_le_n_2);
  gl_gr_lg_le_g368 : AOI21D2BWP7T port map(A1 => CTS_24, A2 => gl_gr_lg_le_n_32, B => gl_gr_lg_le_n_31, ZN => gl_gr_lg_le_n_18);
  gl_gr_lg_le_g369 : CKXOR2D1BWP7T port map(A1 => gl_gr_lg_le_n_32, A2 => gl_sig_e(0), Z => gl_gr_lg_le_n_1);
  gl_gr_lg_le_g370 : ND2D1BWP7T port map(A1 => gl_gr_lg_le_n_32, A2 => gl_sig_e(0), ZN => gl_gr_lg_le_n_0);
  gl_gr_lg_le_count_e_reg_5 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => FE_PHN42_gl_gr_lg_le_new_count_e_5, Q => gl_sig_e(5));
  gl_gr_lg_le_count_e_reg_4 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => FE_PHN46_gl_gr_lg_le_new_count_e_4, Q => gl_sig_e(4));
  gl_gr_lg_le_count_e_reg_0 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => gl_gr_lg_le_new_count_e(0), Q => gl_sig_e(0));
  gl_gr_lg_le_count_e_reg_6 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => FE_PHN41_gl_gr_lg_le_new_count_e_6, Q => gl_sig_e(6));
  gl_gr_lg_le_count_e_reg_7 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => FE_PHN48_gl_gr_lg_le_new_count_e_7, Q => gl_sig_e(7));
  gl_gr_lg_le_count_e_reg_1 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => gl_gr_lg_le_new_count_e(1), Q => gl_sig_e(1));
  gl_gr_lg_le_count_e_reg_9 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => FE_PHN45_gl_gr_lg_le_new_count_e_9, Q => gl_sig_e(9));
  gl_gr_lg_le_count_e_reg_8 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => FE_PHN43_gl_gr_lg_le_new_count_e_8, Q => gl_sig_e(8));
  gl_gr_lg_le_count_e_reg_2 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => FE_PHN47_gl_gr_lg_le_new_count_e_2, Q => gl_sig_e(2));
  gl_gr_lg_le_count_e_reg_3 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => FE_PHN44_gl_gr_lg_le_new_count_e_3, Q => gl_sig_e(3));
  gl_vga_buf_B2_Q_reg : EDFQD0BWP7T port map(CP => CTS_20, D => FE_PHN81_gl_vga_buf_Bint, E => FE_DBTN0_reset, Q => FE_OFN33_B);
  gl_gr_lg_lh_count_h_reg_3 : DFQD0BWP7T port map(CP => CTS_19, D => FE_PHN181_gl_gr_lg_lh_n_17, Q => gl_gr_lg_local_x(3));
  gl_gr_lg_lh_g403 : OAI31D0BWP7T port map(A1 => gl_gr_lg_lh_n_5, A2 => gl_gr_lg_lh_n_3, A3 => gl_gr_lg_lh_n_8, B => gl_gr_lg_lh_n_16, ZN => gl_gr_lg_lh_n_17);
  gl_gr_lg_lh_g405 : OAI21D0BWP7T port map(A1 => gl_gr_lg_lh_n_12, A2 => gl_gr_lg_lh_n_7, B => gl_gr_lg_local_x(3), ZN => gl_gr_lg_lh_n_16);
  gl_gr_lg_lh_g406 : OAI32D0BWP7T port map(A1 => gl_gr_lg_local_x(2), A2 => gl_gr_lg_lh_n_5, A3 => gl_gr_lg_lh_n_8, B1 => gl_gr_lg_lh_n_3, B2 => gl_gr_lg_lh_n_13, ZN => gl_gr_lg_lh_n_15);
  gl_gr_lg_lh_g407 : OAI22D0BWP7T port map(A1 => gl_gr_lg_lh_n_10, A2 => gl_gr_lg_lh_n_5, B1 => gl_gr_lg_lh_n_8, B2 => gl_gr_lg_local_x(1), ZN => gl_gr_lg_lh_n_14);
  gl_gr_lg_lh_g409 : INVD0BWP7T port map(I => gl_gr_lg_lh_n_12, ZN => gl_gr_lg_lh_n_13);
  gl_gr_lg_lh_g410 : IOA21D1BWP7T port map(A1 => gl_gr_lg_lh_n_7, A2 => gl_gr_lg_lh_n_5, B => gl_gr_lg_lh_n_10, ZN => gl_gr_lg_lh_n_12);
  gl_gr_lg_lh_g412 : AOI21D0BWP7T port map(A1 => gl_gr_lg_lh_n_7, A2 => gl_gr_lg_lh_n_4, B => gl_gr_lg_lh_n_6, ZN => gl_gr_lg_lh_n_10);
  gl_gr_lg_lh_g414 : ND3D0BWP7T port map(A1 => gl_gr_lg_lh_n_7, A2 => gl_gr_lg_lh_sig_edges, A3 => gl_gr_lg_local_x(0), ZN => gl_gr_lg_lh_n_8);
  gl_gr_lg_lh_g415 : AOI31D0BWP7T port map(A1 => gl_gr_lg_local_x(2), A2 => gl_gr_lg_local_x(3), A3 => gl_gr_lg_local_x(1), B => FE_OFN35_reset, ZN => gl_gr_lg_lh_n_7);
  gl_gr_lg_lh_g416 : NR2D1BWP7T port map(A1 => gl_gr_lg_lh_sig_edges, A2 => FE_OFN35_reset, ZN => gl_gr_lg_lh_n_6);
  gl_gr_lg_lh_count_h_reg_0 : DFD1BWP7T port map(CP => CTS_19, D => FE_PHN301_gl_gr_lg_lh_n_21, Q => gl_gr_lg_local_x(0), QN => gl_gr_lg_lh_n_4);
  gl_gr_lg_lh_g2 : AO32D1BWP7T port map(A1 => gl_gr_lg_lh_n_7, A2 => gl_gr_lg_lh_sig_edges, A3 => gl_gr_lg_lh_n_4, B1 => gl_gr_lg_lh_n_6, B2 => gl_gr_lg_local_x(0), Z => gl_gr_lg_lh_n_21);
  gl_gr_lg_lh_count_h_reg_1 : DFD1BWP7T port map(CP => CTS_19, D => FE_PHN300_gl_gr_lg_lh_n_14, Q => gl_gr_lg_local_x(1), QN => gl_gr_lg_lh_n_5);
  gl_gr_lg_lh_count_h_reg_2 : DFD1BWP7T port map(CP => CTS_19, D => FE_PHN93_gl_gr_lg_lh_n_15, Q => gl_gr_lg_local_x(2), QN => gl_gr_lg_lh_n_3);
  ml_ms_g754 : OR2D1BWP7T port map(A1 => ml_ms_n_62, A2 => ml_ms_n_63, Z => FE_OFN36_clk15k_switch);
  ml_ms_g755 : INR2XD0BWP7T port map(A1 => ml_ms_sfsm_n_383, B1 => FE_PHN526_ml_ms_muxFSM, ZN => ml_ms_n_63);
  ml_ms_g757 : NR2XD0BWP7T port map(A1 => ml_ms_n_61, A2 => ml_ms_sfsm_state(0), ZN => ml_ms_n_62);
  ml_ms_g758 : CKAN2D1BWP7T port map(A1 => ml_ms_sfsm_state(1), A2 => FE_PHN515_ml_ms_sfsm_state_0, Z => ml_ms_sfsm_n_383);
  ml_ms_g760 : IND2D1BWP7T port map(A1 => ml_ms_sfsm_state(1), B1 => FE_PHN526_ml_ms_muxFSM, ZN => ml_ms_n_61);
  ml_ms_g2 : INR2D1BWP7T port map(A1 => ml_ms_n_61, B1 => ml_ms_sfsm_state(0), ZN => ml_ms_cntReset25M_send);
  ml_ms_sfsm_state_reg_0 : DFQD1BWP7T port map(CP => CTS_20, D => FE_PHN546_ml_ms_n_58, Q => ml_ms_sfsm_state(0));
  ml_ms_sr_new_new_data_reg_0 : DFQD1BWP7T port map(CP => CTS_20, D => FE_PHN548_ml_ms_n_30, Q => ml_ms_sr_new_new_data(0));
  ml_ms_sr_new_new_data_reg_1 : DFQD1BWP7T port map(CP => CTS_20, D => ml_ms_n_20, Q => ml_ms_sr_new_new_data(1));
  ml_ms_sr_new_new_data_reg_2 : DFQD1BWP7T port map(CP => CTS_20, D => ml_ms_n_19, Q => ml_ms_sr_new_new_data(2));
  ml_ms_sr_new_new_data_reg_3 : DFQD1BWP7T port map(CP => CTS_20, D => ml_ms_n_26, Q => ml_ms_sr_new_new_data(3));
  ml_ms_sr_new_new_data_reg_4 : DFQD1BWP7T port map(CP => CTS_20, D => ml_ms_n_25, Q => ml_ms_sr_new_new_data(4));
  ml_ms_sr_new_new_data_reg_5 : DFQD1BWP7T port map(CP => CTS_20, D => FE_PHN550_ml_ms_n_34, Q => ml_ms_sr_new_new_data(5));
  ml_ms_sr_new_new_data_reg_6 : DFQD1BWP7T port map(CP => CTS_20, D => FE_PHN619_ml_ms_n_24, Q => FE_PHN552_ml_ms_sr_new_new_data_6);
  ml_ms_sr_new_new_data_reg_7 : DFQD1BWP7T port map(CP => CTS_20, D => FE_PHN549_ml_ms_n_32, Q => ml_ms_sr_new_new_data(7));
  ml_ms_sr_new_new_data_reg_8 : DFQD1BWP7T port map(CP => CTS_20, D => FE_PHN460_ml_ms_n_31, Q => ml_ms_muxReg);
  ml_ms_g1847 : MOAI22D0BWP7T port map(A1 => ml_ms_n_45, A2 => ml_ms_n_10, B1 => ml_ms_n_59, B2 => FE_PHN446_ml_ms_mux_select, ZN => ml_ms_n_60);
  ml_ms_g1850 : OAI211D1BWP7T port map(A1 => ml_ms_n_8, A2 => ml_ms_n_47, B => ml_ms_n_55, C => ml_ms_n_52, ZN => ml_ms_n_59);
  ml_ms_g1851 : OAI211D1BWP7T port map(A1 => ml_ms_n_49, A2 => ml_ms_n_53, B => ml_ms_n_56, C => ml_ms_n_52, ZN => FE_PHN457_ml_ms_n_58);
  ml_ms_g1852 : OAI221D0BWP7T port map(A1 => ml_ms_n_53, A2 => ml_ms_n_50, B1 => ml_ms_n_0, B2 => ml_ms_n_8, C => ml_ms_n_51, ZN => ml_ms_n_57);
  ml_ms_g1854 : OAI21D0BWP7T port map(A1 => ml_ms_n_47, A2 => ml_ms_n_14, B => ml_ms_n_7, ZN => ml_ms_n_56);
  ml_ms_g1855 : IND3D1BWP7T port map(A1 => ml_ms_n_10, B1 => ml_ms_muxFSM, B2 => ml_ms_n_50, ZN => ml_ms_n_55);
  ml_ms_g1856 : MOAI22D0BWP7T port map(A1 => ml_ms_n_48, A2 => ml_ms_n_16, B1 => ml_ms_n_46, B2 => ml_ms_muxFSM, ZN => FE_PHN379_ml_ms_n_54);
  ml_ms_g1857 : IND3D1BWP7T port map(A1 => ml_ms_n_10, B1 => FE_PHN526_ml_ms_muxFSM, B2 => ml_ms_n_45, ZN => ml_ms_n_53);
  ml_ms_g1858 : IND3D1BWP7T port map(A1 => ml_ms_n_40, B1 => ml_ms_n_45, B2 => ml_ms_n_48, ZN => ml_ms_n_51);
  ml_ms_g1859 : IND3D1BWP7T port map(A1 => ml_ms_n_16, B1 => ml_ms_n_37, B2 => ml_ms_n_48, ZN => ml_ms_n_52);
  ml_ms_g1860 : INVD0BWP7T port map(I => ml_ms_n_50, ZN => ml_ms_n_49);
  ml_ms_g1861 : IAO21D0BWP7T port map(A1 => ml_ms_n_43, A2 => ml_ms_n_11, B => ml_ms_count25M(12), ZN => ml_ms_n_50);
  ml_ms_g1862 : IOA21D1BWP7T port map(A1 => ml_ms_n_42, A2 => ml_ms_n_18, B => ml_ms_sfsm_state(1), ZN => ml_ms_n_48);
  ml_ms_g1863 : AOI21D0BWP7T port map(A1 => ml_ms_n_44, A2 => ml_ms_sfsm_state(0), B => ml_ms_reset_send, ZN => ml_ms_n_46);
  ml_ms_g1864 : AOI211XD0BWP7T port map(A1 => ml_ms_sfsm_state(1), A2 => clk15k_in, B => ml_ms_n_41, C => ml_ms_n_1, ZN => ml_ms_n_47);
  ml_ms_g1865 : ND2D1BWP7T port map(A1 => ml_ms_n_44, A2 => FE_PHN526_ml_ms_muxFSM, ZN => ml_ms_n_45);
  ml_ms_g1866 : NR2XD0BWP7T port map(A1 => ml_ms_n_38, A2 => FE_PHN323_ml_ms_count25M_9, ZN => ml_ms_n_43);
  ml_ms_g1867 : OA31D1BWP7T port map(A1 => ml_ms_count25M(11), A2 => ml_ms_count25M(10), A3 => ml_ms_n_33, B => ml_ms_sfsm_state(1), Z => ml_ms_n_44);
  ml_ms_g1868 : OAI211D1BWP7T port map(A1 => ml_ms_n_17, A2 => ml_ms_n_36, B => ml_ms_count25M(11), C => FE_PHN323_ml_ms_count25M_9, ZN => ml_ms_n_42);
  ml_ms_g1869 : NR2D1BWP7T port map(A1 => ml_ms_n_39, A2 => ml_ms_sfsm_state(1), ZN => ml_ms_n_41);
  ml_ms_g1870 : OA22D0BWP7T port map(A1 => ml_ms_n_16, A2 => ml_ms_n_37, B1 => ml_ms_n_0, B2 => ml_ms_n_10, Z => ml_ms_n_40);
  ml_ms_g1871 : AOI21D0BWP7T port map(A1 => ml_ms_n_35, A2 => ml_ms_n_15, B => ml_ms_n_18, ZN => ml_ms_n_39);
  ml_ms_g1872 : AO211D0BWP7T port map(A1 => ml_ms_n_27, A2 => ml_ms_count25M(8), B => ml_ms_n_29, C => ml_ms_n_17, Z => ml_ms_n_38);
  ml_ms_g1877 : ND4D0BWP7T port map(A1 => ml_ms_n_12, A2 => ml_ms_count25M(8), A3 => FE_PHN323_ml_ms_count25M_9, A4 => ml_ms_count25M(12), ZN => ml_ms_n_37);
  ml_ms_g1878 : AN2D0BWP7T port map(A1 => ml_ms_n_29, A2 => ml_ms_count25M(3), Z => ml_ms_n_36);
  ml_ms_g1884 : OAI211D1BWP7T port map(A1 => ml_ms_count25M(3), A2 => ml_ms_n_3, B => ml_ms_n_5, C => ml_ms_count25M(5), ZN => ml_ms_n_35);
  ml_ms_g1885 : ND2D1BWP7T port map(A1 => ml_ms_n_28, A2 => FE_PHN618_ml_ms_n_22, ZN => ml_ms_n_34);
  ml_ms_g1886 : OAI21D0BWP7T port map(A1 => ml_ms_n_13, A2 => ml_ms_n_6, B => ml_ms_n_15, ZN => ml_ms_n_33);
  ml_ms_g1887 : ND2D1BWP7T port map(A1 => ml_ms_n_28, A2 => ml_ms_n_23, ZN => ml_ms_n_32);
  ml_ms_g1888 : ND2D1BWP7T port map(A1 => ml_ms_n_28, A2 => ml_ms_n_21, ZN => ml_ms_n_31);
  ml_ms_g1889 : IOA21D1BWP7T port map(A1 => ml_ms_n_4, A2 => FE_PHN623_ml_ms_sr_new_new_data_0, B => ml_ms_n_28, ZN => ml_ms_n_30);
  ml_ms_g1890 : AN4D0BWP7T port map(A1 => ml_ms_count25M(3), A2 => ml_ms_count25M(2), A3 => ml_ms_count25M(7), A4 => ml_ms_count25M(5), Z => ml_ms_n_27);
  ml_ms_g1891 : AO22D0BWP7T port map(A1 => ml_ms_n_4, A2 => ml_ms_sr_new_new_data(3), B1 => ml_ms_sr_new_new_data(2), B2 => ml_ms_n_9, Z => FE_PHN77_ml_ms_n_26);
  ml_ms_g1892 : AO22D0BWP7T port map(A1 => ml_ms_n_4, A2 => ml_ms_sr_new_new_data(4), B1 => ml_ms_sr_new_new_data(3), B2 => ml_ms_n_9, Z => FE_PHN73_ml_ms_n_25);
  ml_ms_g1893 : AN4D0BWP7T port map(A1 => ml_ms_count25M(4), A2 => ml_ms_count25M(8), A3 => ml_ms_count25M(7), A4 => ml_ms_count25M(5), Z => ml_ms_n_29);
  ml_ms_g1894 : OAI211D1BWP7T port map(A1 => FE_PHN526_ml_ms_muxFSM, A2 => ml_ms_sfsm_n_383, B => ml_ms_actBit, C => FE_PHN441_ml_ms_n_2, ZN => ml_ms_n_28);
  ml_ms_g1895 : AO22D0BWP7T port map(A1 => ml_ms_n_4, A2 => ml_ms_sr_new_new_data(6), B1 => FE_PHN516_ml_ms_sr_new_new_data_5, B2 => ml_ms_n_9, Z => ml_ms_n_24);
  ml_ms_g1896 : AOI22D0BWP7T port map(A1 => ml_ms_n_4, A2 => FE_PHN466_ml_ms_sr_new_new_data_7, B1 => ml_ms_n_9, B2 => ml_ms_sr_new_new_data(6), ZN => FE_PHN620_ml_ms_n_23);
  ml_ms_g1897 : AOI22D0BWP7T port map(A1 => ml_ms_n_4, A2 => FE_PHN516_ml_ms_sr_new_new_data_5, B1 => ml_ms_n_9, B2 => FE_PHN641_ml_ms_sr_new_new_data_4, ZN => ml_ms_n_22);
  ml_ms_g1898 : AOI22D0BWP7T port map(A1 => ml_ms_n_4, A2 => FE_PHN566_ml_ms_muxReg, B1 => ml_ms_n_9, B2 => FE_PHN466_ml_ms_sr_new_new_data_7, ZN => FE_PHN545_ml_ms_n_21);
  ml_ms_g1899 : AO22D0BWP7T port map(A1 => ml_ms_n_4, A2 => ml_ms_sr_new_new_data(1), B1 => ml_ms_sr_new_new_data(0), B2 => ml_ms_n_9, Z => FE_PHN75_ml_ms_n_20);
  ml_ms_g1900 : AO22D0BWP7T port map(A1 => ml_ms_n_4, A2 => ml_ms_sr_new_new_data(2), B1 => ml_ms_sr_new_new_data(1), B2 => ml_ms_n_9, Z => FE_PHN74_ml_ms_n_19);
  ml_ms_g1901 : INR2D1BWP7T port map(A1 => ml_ms_n_11, B1 => ml_ms_count25M(12), ZN => ml_ms_n_18);
  ml_ms_g1902 : INR2D1BWP7T port map(A1 => ml_ms_count25M(8), B1 => ml_ms_n_6, ZN => ml_ms_n_17);
  ml_ms_g1903 : OR2D1BWP7T port map(A1 => ml_ms_n_10, A2 => ml_ms_muxFSM, Z => ml_ms_n_16);
  ml_ms_g1904 : AOI21D0BWP7T port map(A1 => ml_ms_n_0, A2 => FE_PHN446_ml_ms_mux_select, B => FE_PHN526_ml_ms_muxFSM, ZN => ml_ms_n_14);
  ml_ms_g1905 : NR3D0BWP7T port map(A1 => ml_ms_count25M(3), A2 => ml_ms_count25M(4), A3 => ml_ms_count25M(5), ZN => ml_ms_n_13);
  ml_ms_g1906 : IAO21D0BWP7T port map(A1 => ml_ms_count25M(7), A2 => FE_PHN318_ml_ms_count25M_6, B => ml_ms_n_11, ZN => ml_ms_n_12);
  ml_ms_g1907 : NR3D0BWP7T port map(A1 => ml_ms_count25M(8), A2 => ml_ms_count25M(12), A3 => FE_PHN323_ml_ms_count25M_9, ZN => ml_ms_n_15);
  ml_ms_g1908 : ND2D1BWP7T port map(A1 => ml_ms_count25M(10), A2 => ml_ms_count25M(11), ZN => ml_ms_n_11);
  ml_ms_g1909 : IND2D1BWP7T port map(A1 => ml_ms_reset_send, B1 => FE_PHN515_ml_ms_sfsm_state_0, ZN => ml_ms_n_10);
  ml_ms_g1910 : AN2D1BWP7T port map(A1 => ml_ms_output_edgedet, A2 => FE_PHN446_ml_ms_mux_select, Z => ml_ms_n_9);
  ml_ms_g1911 : INVD1BWP7T port map(I => ml_ms_n_7, ZN => ml_ms_n_8);
  ml_ms_g1912 : INVD0BWP7T port map(I => ml_ms_n_6, ZN => ml_ms_n_5);
  ml_ms_g1913 : OR2D1BWP7T port map(A1 => ml_ms_count25M(4), A2 => ml_ms_count25M(2), Z => ml_ms_n_3);
  ml_ms_g1914 : NR2XD0BWP7T port map(A1 => ml_ms_reset_send, A2 => ml_ms_sfsm_state(0), ZN => ml_ms_n_7);
  ml_ms_g1915 : CKND2D1BWP7T port map(A1 => ml_ms_count25M(7), A2 => FE_PHN318_ml_ms_count25M_6, ZN => ml_ms_n_6);
  ml_ms_g1916 : NR2XD0BWP7T port map(A1 => ml_ms_output_edgedet, A2 => FE_PHN441_ml_ms_n_2, ZN => ml_ms_n_4);
  ml_ms_sfsm_state_reg_1 : DFD1BWP7T port map(CP => CTS_20, D => FE_PHN372_ml_ms_n_57, Q => ml_ms_sfsm_state(1), QN => ml_ms_n_0);
  ml_ms_sfsm_state_reg_3 : DFD1BWP7T port map(CP => CTS_20, D => FE_PHN544_ml_ms_n_60, Q => ml_ms_mux_select, QN => ml_ms_n_2);
  ml_ms_sfsm_state_reg_2 : DFD1BWP7T port map(CP => CTS_20, D => ml_ms_n_54, Q => ml_ms_muxFSM, QN => ml_ms_n_1);
  ml_ms_mfsm_g2156 : IND4D0BWP7T port map(A1 => ml_ms_mfsm_n_118, B1 => ml_ms_mfsm_n_56, B2 => ml_ms_mfsm_n_62, B3 => ml_ms_mfsm_n_63, ZN => ml_ms_cntReset15K);
  ml_ms_mfsm_g2157 : AN2D0BWP7T port map(A1 => ml_ms_btnflipfloprst, A2 => ml_ms_data_sr_11bit(3), Z => ml_ms_btns(4));
  ml_ms_mfsm_g2158 : AN2D0BWP7T port map(A1 => ml_ms_btnflipfloprst, A2 => ml_ms_data_sr_11bit(4), Z => ml_ms_btns(3));
  ml_ms_mfsm_g2159 : AN2D0BWP7T port map(A1 => ml_ms_btnflipfloprst, A2 => FE_PHN279_ml_ms_data_sr_11bit_2, Z => ml_ms_btns(2));
  ml_ms_mfsm_g2160 : AN2D0BWP7T port map(A1 => ml_ms_btnflipfloprst, A2 => ml_ms_data_sr_11bit(7), Z => ml_ms_btns(1));
  ml_ms_mfsm_g2161 : AN2D0BWP7T port map(A1 => ml_ms_btnflipfloprst, A2 => ml_ms_data_sr_11bit(6), Z => ml_ms_btns(0));
  ml_ms_mfsm_g2162 : INR2D1BWP7T port map(A1 => FE_PHN279_ml_ms_data_sr_11bit_2, B1 => ml_ms_mfsm_n_64, ZN => ml_ms_mouse_x(0));
  ml_ms_mfsm_g2163 : INR2D1BWP7T port map(A1 => ml_ms_data_sr_11bit(3), B1 => ml_ms_mfsm_n_64, ZN => ml_ms_mouse_x(1));
  ml_ms_mfsm_g2164 : INR2D1BWP7T port map(A1 => ml_ms_data_sr_11bit(4), B1 => ml_ms_mfsm_n_64, ZN => ml_ms_mouse_x(2));
  ml_ms_mfsm_g2165 : AN2D0BWP7T port map(A1 => ml_ms_yflipfloprst, A2 => ml_ms_data_sr_11bit(4), Z => ml_ms_mouse_y(2));
  ml_ms_mfsm_g2166 : AN2D0BWP7T port map(A1 => ml_ms_yflipfloprst, A2 => ml_ms_data_sr_11bit(3), Z => ml_ms_mouse_y(1));
  ml_ms_mfsm_g2167 : AN2D0BWP7T port map(A1 => ml_ms_yflipfloprst, A2 => FE_PHN279_ml_ms_data_sr_11bit_2, Z => ml_ms_mouse_y(0));
  ml_ms_mfsm_g2168 : ND3D0BWP7T port map(A1 => ml_ms_mfsm_n_61, A2 => ml_ms_mfsm_n_60, A3 => ml_ms_mfsm_state(1), ZN => ml_ms_cntReset25M_main);
  ml_ms_mfsm_g2169 : OAI31D1BWP7T port map(A1 => FE_PHN338_ml_ms_mfsm_state_2, A2 => FE_PHN347_ml_ms_mfsm_state_3, A3 => ml_ms_mfsm_n_59, B => ml_ms_mfsm_n_62, ZN => ml_ms_btnflipfloprst);
  ml_ms_mfsm_g2170 : NR2XD0BWP7T port map(A1 => ml_ms_reset_send, A2 => ml_ms_mfsm_n_1, ZN => ml_ms_actBit);
  ml_ms_mfsm_g2171 : IAO21D0BWP7T port map(A1 => ml_ms_mfsm_n_59, A2 => ml_ms_mfsm_n_53, B => ml_ms_xflipfloprst, ZN => ml_ms_mfsm_n_64);
  ml_ms_mfsm_g2172 : AO211D0BWP7T port map(A1 => ml_ms_mfsm_n_57, A2 => ml_ms_mfsm_n_3, B => ml_ms_mfsm_n_55, C => ml_ms_mfsm_n_54, Z => ml_ms_mux_select_main);
  ml_ms_mfsm_g2173 : AOI22D0BWP7T port map(A1 => ml_ms_mfsm_n_58, A2 => FE_PHN347_ml_ms_mfsm_state_3, B1 => ml_ms_mfsm_n_55, B2 => ml_ms_mfsm_n_4, ZN => ml_ms_mfsm_n_63);
  ml_ms_mfsm_g2174 : MOAI22D0BWP7T port map(A1 => ml_ms_mfsm_n_117, A2 => ml_ms_mfsm_n_56, B1 => ml_ms_mfsm_n_118, B2 => FE_PHN338_ml_ms_mfsm_state_2, ZN => ml_ms_yflipfloprst);
  ml_ms_mfsm_g2175 : AN2D1BWP7T port map(A1 => ml_ms_mfsm_n_118, A2 => FE_PHN329_ml_ms_mfsm_n_53, Z => ml_ms_xflipfloprst);
  ml_ms_mfsm_g2176 : ND2D1BWP7T port map(A1 => ml_ms_mfsm_n_116, A2 => FE_PHN338_ml_ms_mfsm_state_2, ZN => ml_ms_mfsm_n_62);
  ml_ms_mfsm_g2177 : AOI22D0BWP7T port map(A1 => ml_ms_mfsm_n_55, A2 => ml_ms_mfsm_state(2), B1 => ml_ms_mfsm_n_53, B2 => ml_ms_mfsm_state(3), ZN => ml_ms_mfsm_n_61);
  ml_ms_mfsm_g2178 : MAOI22D0BWP7T port map(A1 => ml_ms_mfsm_n_54, A2 => ml_ms_mfsm_n_4, B1 => ml_ms_mfsm_n_54, B2 => ml_ms_mfsm_n_4, ZN => ml_ms_mfsm_n_60);
  ml_ms_mfsm_g2179 : ND3D0BWP7T port map(A1 => ml_ms_mfsm_n_54, A2 => ml_ms_mfsm_n_0, A3 => ml_ms_mfsm_state(0), ZN => ml_ms_reset_send);
  ml_ms_mfsm_g2180 : ND2D1BWP7T port map(A1 => ml_ms_mfsm_n_57, A2 => FE_PHN350_ml_ms_mfsm_state_4, ZN => ml_ms_mfsm_n_59);
  ml_ms_mfsm_g2181 : AN2D1BWP7T port map(A1 => ml_ms_mfsm_n_66, A2 => FE_PHN350_ml_ms_mfsm_state_4, Z => ml_ms_mfsm_n_118);
  ml_ms_mfsm_g2182 : NR2XD0BWP7T port map(A1 => ml_ms_mfsm_n_56, A2 => ml_ms_mfsm_n_4, ZN => ml_handshake_mouse_out);
  ml_ms_mfsm_g2183 : OAI21D0BWP7T port map(A1 => ml_ms_mfsm_state(0), A2 => FE_PHN338_ml_ms_mfsm_state_2, B => ml_ms_mfsm_n_117, ZN => ml_ms_mfsm_n_58);
  ml_ms_mfsm_g2184 : AN2D1BWP7T port map(A1 => ml_ms_mfsm_n_66, A2 => FE_PHN347_ml_ms_mfsm_state_3, Z => ml_ms_mfsm_n_116);
  ml_ms_mfsm_g2185 : INVD0BWP7T port map(I => ml_ms_mfsm_n_57, ZN => ml_ms_mfsm_n_117);
  ml_ms_mfsm_g2186 : NR2XD0BWP7T port map(A1 => ml_ms_mfsm_n_0, A2 => ml_ms_mfsm_n_4, ZN => ml_ms_mfsm_n_66);
  ml_ms_mfsm_g2187 : NR2XD0BWP7T port map(A1 => ml_ms_mfsm_state(1), A2 => ml_ms_mfsm_state(0), ZN => ml_ms_mfsm_n_57);
  ml_ms_mfsm_g2188 : ND2D1BWP7T port map(A1 => FE_PHN347_ml_ms_mfsm_state_3, A2 => FE_PHN350_ml_ms_mfsm_state_4, ZN => ml_ms_mfsm_n_56);
  ml_ms_mfsm_g2189 : NR2D0BWP7T port map(A1 => ml_ms_mfsm_state(3), A2 => FE_PHN350_ml_ms_mfsm_state_4, ZN => ml_ms_mfsm_n_55);
  ml_ms_mfsm_g2190 : NR2XD0BWP7T port map(A1 => ml_ms_mfsm_state(2), A2 => FE_PHN350_ml_ms_mfsm_state_4, ZN => ml_ms_mfsm_n_54);
  ml_ms_mfsm_g2722 : OAI21D0BWP7T port map(A1 => ml_ms_mfsm_n_33, A2 => FE_PHN350_ml_ms_mfsm_state_4, B => ml_ms_mfsm_n_51, ZN => ml_ms_mfsm_n_52);
  ml_ms_mfsm_g2723 : AOI22D0BWP7T port map(A1 => ml_ms_mfsm_n_49, A2 => ml_ms_mfsm_n_8, B1 => ml_ms_mfsm_n_50, B2 => ml_ms_mfsm_n_17, ZN => ml_ms_mfsm_n_51);
  ml_ms_mfsm_g2724 : AOI211XD0BWP7T port map(A1 => ml_ms_mfsm_n_14, A2 => ml_ms_mfsm_n_4, B => ml_ms_mfsm_n_48, C => ml_ms_mfsm_n_29, ZN => ml_ms_mfsm_n_50);
  ml_ms_mfsm_g2725 : OAI22D0BWP7T port map(A1 => ml_ms_mfsm_n_47, A2 => FE_PHN350_ml_ms_mfsm_state_4, B1 => ml_ms_mfsm_n_45, B2 => ml_ms_mfsm_n_14, ZN => ml_ms_mfsm_n_49);
  ml_ms_mfsm_g2726 : OAI32D1BWP7T port map(A1 => ml_ms_mfsm_state(1), A2 => ml_ms_mfsm_n_4, A3 => ml_ms_mfsm_n_10, B1 => FE_PHN347_ml_ms_mfsm_state_3, B2 => ml_ms_mfsm_n_46, ZN => ml_ms_mfsm_n_48);
  ml_ms_mfsm_g2728 : AOI22D0BWP7T port map(A1 => ml_ms_mfsm_n_43, A2 => FE_PHN347_ml_ms_mfsm_state_3, B1 => ml_ms_mfsm_n_28, B2 => ml_ms_mfsm_n_1, ZN => ml_ms_mfsm_n_47);
  ml_ms_mfsm_g2730 : INVD0BWP7T port map(I => ml_ms_mfsm_n_45, ZN => ml_ms_mfsm_n_46);
  ml_ms_mfsm_g2731 : OAI31D0BWP7T port map(A1 => ml_ms_mfsm_n_4, A2 => ml_ms_mfsm_n_10, A3 => ml_ms_mfsm_n_18, B => ml_ms_mfsm_n_41, ZN => ml_ms_mfsm_n_44);
  ml_ms_mfsm_g2732 : ND2D1BWP7T port map(A1 => ml_ms_mfsm_n_43, A2 => ml_ms_mfsm_n_28, ZN => ml_ms_mfsm_n_45);
  ml_ms_mfsm_g2733 : AOI31D0BWP7T port map(A1 => ml_ms_mfsm_n_34, A2 => ml_ms_mfsm_n_5, A3 => ml_ms_mfsm_state(1), B => ml_ms_mfsm_n_66, ZN => ml_ms_mfsm_n_43);
  ml_ms_mfsm_g2735 : OAI211D1BWP7T port map(A1 => FE_PHN320_ml_buttons_mouse_3, A2 => ml_ms_mfsm_n_26, B => ml_ms_mfsm_n_39, C => ml_ms_mfsm_n_22, ZN => ml_ms_mfsm_n_42);
  ml_ms_mfsm_g2736 : AOI31D0BWP7T port map(A1 => ml_ms_mfsm_n_32, A2 => ml_ms_mfsm_n_6, A3 => ml_ms_mfsm_n_3, B => ml_ms_mfsm_n_40, ZN => ml_ms_mfsm_n_41);
  ml_ms_mfsm_g2737 : AO222D0BWP7T port map(A1 => ml_ms_mfsm_n_31, A2 => ml_ms_mfsm_n_23, B1 => ml_ms_mfsm_n_15, B2 => ml_ms_mfsm_n_17, C1 => ml_ms_mfsm_n_30, C2 => ml_ms_mfsm_n_25, Z => ml_ms_mfsm_n_40);
  ml_ms_mfsm_g2738 : AOI211XD0BWP7T port map(A1 => ml_ms_mfsm_n_29, A2 => ml_ms_mfsm_n_6, B => ml_ms_mfsm_n_37, C => ml_ms_mfsm_n_19, ZN => ml_ms_mfsm_n_39);
  ml_ms_mfsm_g2739 : OAI22D0BWP7T port map(A1 => ml_ms_mfsm_n_35, A2 => ml_ms_mfsm_n_9, B1 => ml_ms_mfsm_n_13, B2 => ml_ms_mfsm_n_1, ZN => ml_ms_mfsm_n_38);
  ml_ms_mfsm_g2741 : NR4D0BWP7T port map(A1 => ml_ms_mfsm_n_29, A2 => ml_ms_mfsm_n_116, A3 => ml_ms_mfsm_n_9, A4 => FE_PHN350_ml_ms_mfsm_state_4, ZN => ml_ms_mfsm_n_37);
  ml_ms_mfsm_g2742 : OAI211D1BWP7T port map(A1 => ml_ms_mfsm_n_3, A2 => ml_ms_mfsm_n_27, B => ml_ms_mfsm_n_16, C => ml_ms_mfsm_n_18, ZN => ml_ms_mfsm_n_36);
  ml_ms_mfsm_g2743 : AOI21D0BWP7T port map(A1 => ml_ms_mfsm_n_29, A2 => ml_ms_mfsm_n_1, B => ml_ms_mfsm_n_118, ZN => ml_ms_mfsm_n_35);
  ml_ms_mfsm_g2744 : OAI31D0BWP7T port map(A1 => FE_PHN323_ml_ms_count25M_9, A2 => ml_ms_count25M(10), A3 => ml_ms_mfsm_n_24, B => ml_ms_count25M(11), ZN => ml_ms_mfsm_n_34);
  ml_ms_mfsm_g2745 : IND3D1BWP7T port map(A1 => ml_ms_mfsm_n_29, B1 => ml_ms_mfsm_n_6, B2 => FE_PHN467_ml_ms_mfsm_n_21, ZN => ml_ms_mfsm_n_33);
  ml_ms_mfsm_g2746 : IOA21D1BWP7T port map(A1 => ml_ms_mfsm_n_28, A2 => ml_ms_mfsm_state(1), B => ml_ms_mfsm_n_21, ZN => ml_ms_mfsm_n_32);
  ml_ms_mfsm_g2747 : OAI21D0BWP7T port map(A1 => ml_ms_mfsm_n_26, A2 => ml_ms_mfsm_n_4, B => ml_ms_mfsm_n_20, ZN => ml_ms_mfsm_n_31);
  ml_ms_mfsm_g2748 : MOAI22D0BWP7T port map(A1 => ml_ms_mfsm_n_28, A2 => ml_ms_mfsm_state(1), B1 => ml_ms_mfsm_n_4, B2 => ml_ms_mfsm_state(1), ZN => ml_ms_mfsm_n_30);
  ml_ms_mfsm_g2749 : NR2XD0BWP7T port map(A1 => ml_ms_mfsm_n_28, A2 => FE_PHN454_ml_ms_mfsm_n_0, ZN => ml_ms_mfsm_n_29);
  ml_ms_mfsm_g2750 : OAI31D0BWP7T port map(A1 => ml_ms_mfsm_state(0), A2 => ml_ms_mfsm_n_0, A3 => ml_ms_mfsm_n_7, B => FE_DBTN0_reset, ZN => ml_ms_mfsm_n_27);
  ml_ms_mfsm_g2751 : OR2D1BWP7T port map(A1 => ml_ms_mfsm_n_23, A2 => ml_ms_mfsm_n_4, Z => ml_ms_mfsm_n_28);
  ml_ms_mfsm_g2752 : IOA21D1BWP7T port map(A1 => ml_ms_mfsm_n_17, A2 => ml_ms_mfsm_n_1, B => ml_ms_mfsm_n_9, ZN => ml_ms_mfsm_n_25);
  ml_ms_mfsm_g2753 : AN4D0BWP7T port map(A1 => ml_ms_mfsm_n_11, A2 => ml_ms_count25M(8), A3 => FE_PHN318_ml_ms_count25M_6, A4 => ml_ms_count25M(7), Z => ml_ms_mfsm_n_24);
  ml_ms_mfsm_g2754 : IND3D1BWP7T port map(A1 => FE_PHN454_ml_ms_mfsm_n_0, B1 => FE_PHN347_ml_ms_mfsm_state_3, B2 => ml_ms_mfsm_n_17, ZN => ml_ms_mfsm_n_26);
  ml_ms_mfsm_g2755 : ND2D1BWP7T port map(A1 => ml_ms_mfsm_n_17, A2 => ml_ms_mfsm_n_66, ZN => ml_ms_mfsm_n_22);
  ml_ms_mfsm_g2756 : IND2D1BWP7T port map(A1 => ml_ms_mfsm_n_12, B1 => ml_ms_count15k(3), ZN => ml_ms_mfsm_n_23);
  ml_ms_mfsm_g2757 : ND4D0BWP7T port map(A1 => ml_ms_mfsm_n_8, A2 => ml_ms_mfsm_n_3, A3 => ml_ms_mfsm_n_1, A4 => ml_ms_mfsm_state(1), ZN => ml_ms_mfsm_n_20);
  ml_ms_mfsm_g2758 : AOI21D0BWP7T port map(A1 => ml_ms_mfsm_n_66, A2 => ml_ms_mfsm_n_7, B => ml_ms_mfsm_n_18, ZN => ml_ms_mfsm_n_19);
  ml_ms_mfsm_g2759 : ND4D0BWP7T port map(A1 => FE_PHN454_ml_ms_mfsm_n_0, A2 => ml_ms_count15k(3), A3 => ml_ms_count15k(2), A4 => ml_ms_mfsm_state(0), ZN => ml_ms_mfsm_n_21);
  ml_ms_mfsm_g2760 : CKND2D0BWP7T port map(A1 => ml_ms_mfsm_n_116, A2 => ml_ms_mfsm_n_8, ZN => ml_ms_mfsm_n_16);
  ml_ms_mfsm_g2761 : INR2D1BWP7T port map(A1 => ml_ms_mfsm_n_117, B1 => ml_ms_mfsm_n_10, ZN => ml_ms_mfsm_n_15);
  ml_ms_mfsm_g2762 : ND2D1BWP7T port map(A1 => ml_ms_mfsm_n_8, A2 => FE_PHN350_ml_ms_mfsm_state_4, ZN => ml_ms_mfsm_n_18);
  ml_ms_mfsm_g2763 : AN2D1BWP7T port map(A1 => ml_ms_mfsm_n_6, A2 => FE_PHN350_ml_ms_mfsm_state_4, Z => ml_ms_mfsm_n_17);
  ml_ms_mfsm_g2764 : IAO21D0BWP7T port map(A1 => ml_ms_mfsm_n_66, A2 => FE_OFN35_reset, B => ml_ms_mfsm_n_6, ZN => ml_ms_mfsm_n_13);
  ml_ms_mfsm_g2765 : AOI21D0BWP7T port map(A1 => ml_ms_count15k(0), A2 => FE_PHN335_ml_ms_count15k_1, B => ml_ms_count15k(2), ZN => ml_ms_mfsm_n_12);
  ml_ms_mfsm_g2766 : OR4D1BWP7T port map(A1 => ml_ms_count25M(5), A2 => ml_ms_count25M(4), A3 => ml_ms_count25M(3), A4 => ml_ms_count25M(2), Z => ml_ms_mfsm_n_11);
  ml_ms_mfsm_g2767 : NR2XD0BWP7T port map(A1 => ml_ms_mfsm_n_10, A2 => FE_PHN454_ml_ms_mfsm_n_0, ZN => ml_ms_mfsm_n_14);
  ml_ms_mfsm_g2768 : INVD1BWP7T port map(I => ml_ms_mfsm_n_9, ZN => ml_ms_mfsm_n_8);
  ml_ms_mfsm_g2769 : ND2D1BWP7T port map(A1 => FE_PHN320_ml_buttons_mouse_3, A2 => FE_PHN347_ml_ms_mfsm_state_3, ZN => ml_ms_mfsm_n_10);
  ml_ms_mfsm_g2770 : ND2D1BWP7T port map(A1 => FE_PHN338_ml_ms_mfsm_state_2, A2 => FE_DBTN0_reset, ZN => ml_ms_mfsm_n_9);
  ml_ms_mfsm_g2771 : OR2D1BWP7T port map(A1 => ml_ms_mfsm_n_1, A2 => FE_PHN320_ml_buttons_mouse_3, Z => ml_ms_mfsm_n_7);
  ml_ms_mfsm_g2772 : NR2D1BWP7T port map(A1 => FE_PHN338_ml_ms_mfsm_state_2, A2 => FE_OFN35_reset, ZN => ml_ms_mfsm_n_6);
  ml_ms_mfsm_g2773 : CKND1BWP7T port map(I => ml_ms_count25M(12), ZN => ml_ms_mfsm_n_5);
  ml_ms_mfsm_state_reg_1 : DFD1BWP7T port map(CP => CTS_20, D => FE_PHN394_ml_ms_mfsm_n_44, Q => ml_ms_mfsm_state(1), QN => ml_ms_mfsm_n_0);
  ml_ms_mfsm_state_reg_0 : DFD1BWP7T port map(CP => CTS_20, D => FE_PHN456_ml_ms_mfsm_n_52, Q => ml_ms_mfsm_state(0), QN => ml_ms_mfsm_n_4);
  ml_ms_mfsm_state_reg_2 : DFD1BWP7T port map(CP => CTS_20, D => ml_ms_mfsm_n_42, Q => ml_ms_mfsm_state(2), QN => ml_ms_mfsm_n_53);
  ml_ms_mfsm_state_reg_4 : DFD1BWP7T port map(CP => CTS_20, D => FE_PHN367_ml_ms_mfsm_n_36, Q => ml_ms_mfsm_state(4), QN => ml_ms_mfsm_n_3);
  ml_ms_mfsm_state_reg_3 : DFD1BWP7T port map(CP => CTS_20, D => FE_PHN387_ml_ms_mfsm_n_38, Q => ml_ms_mfsm_state(3), QN => ml_ms_mfsm_n_1);
  ml_ms_tb_count_reg_3 : EDFKCNQD1BWP7T port map(CN => ml_ms_tb_n_1, CP => CTS_20, D => ml_ms_tb_n_6, E => ml_ms_output_edgedet, Q => ml_ms_count15k(3));
  ml_ms_tb_count_reg_2 : EDFKCNQD1BWP7T port map(CN => ml_ms_tb_n_1, CP => CTS_20, D => ml_ms_tb_n_5, E => ml_ms_output_edgedet, Q => ml_ms_count15k(2));
  ml_ms_tb_g65 : MOAI22D0BWP7T port map(A1 => ml_ms_tb_n_4, A2 => ml_ms_count15k(3), B1 => ml_ms_tb_n_4, B2 => ml_ms_count15k(3), ZN => FE_PHN388_ml_ms_tb_n_6);
  ml_ms_tb_count_reg_1 : EDFKCNQD1BWP7T port map(CN => ml_ms_tb_n_1, CP => CTS_20, D => ml_ms_tb_n_3, E => ml_ms_output_edgedet, Q => ml_ms_count15k(1));
  ml_ms_tb_g67 : MOAI22D0BWP7T port map(A1 => ml_ms_tb_n_2, A2 => ml_ms_count15k(2), B1 => ml_ms_tb_n_2, B2 => ml_ms_count15k(2), ZN => FE_PHN391_ml_ms_tb_n_5);
  ml_ms_tb_count_reg_0 : DFKCNQD1BWP7T port map(CN => ml_ms_tb_n_0, CP => CTS_20, D => ml_ms_tb_n_1, Q => FE_PHN334_ml_ms_count15k_0);
  ml_ms_tb_g69 : IND2D1BWP7T port map(A1 => ml_ms_tb_n_2, B1 => ml_ms_count15k(2), ZN => ml_ms_tb_n_4);
  ml_ms_tb_g70 : CKXOR2D2BWP7T port map(A1 => FE_PHN335_ml_ms_count15k_1, A2 => ml_ms_count15k(0), Z => ml_ms_tb_n_3);
  ml_ms_tb_g72 : ND2D1BWP7T port map(A1 => FE_PHN335_ml_ms_count15k_1, A2 => ml_ms_count15k(0), ZN => ml_ms_tb_n_2);
  ml_ms_tb_g73 : INVD1BWP7T port map(I => ml_ms_cntReset15K, ZN => ml_ms_tb_n_1);
  ml_ms_tb_g2 : CKXOR2D1BWP7T port map(A1 => ml_ms_output_edgedet, A2 => ml_ms_count15k(0), Z => FE_PHN448_ml_ms_tb_n_0);
  ml_ms_flipflop1_Q_reg : DFXQD1BWP7T port map(CP => CTS_19, DA => ml_ms_mouse_x(2), DB => FE_PHN85_ml_mouseX_2, Q => ml_mouseX(2), SA => ml_ms_xflipfloprst);
  ml_ms_flipflop10_Q_reg : EDFQD1BWP7T port map(CP => CTS_20, D => ml_ms_btns(1), E => ml_ms_btnflipfloprst, Q => ml_buttons_mouse(1));
  ml_ms_flipflop2_Q_reg : DFXQD1BWP7T port map(CP => CTS_19, DA => ml_ms_mouse_x(1), DB => FE_PHN84_ml_mouseX_1, Q => ml_mouseX(1), SA => ml_ms_xflipfloprst);
  ml_ms_flipflop11_Q_reg : EDFQD1BWP7T port map(CP => CTS_20, D => ml_ms_btns(0), E => ml_ms_btnflipfloprst, Q => ml_buttons_mouse(0));
  ml_ms_flipflop3_Q_reg : DFXQD1BWP7T port map(CP => CTS_20, DA => ml_ms_mouse_x(0), DB => FE_PHN76_ml_mouseX_0, Q => ml_mouseX(0), SA => ml_ms_xflipfloprst);
  ml_ms_sr11_data_out_reg_1 : EDFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_20, D => FE_PHN86_ml_ms_sr11_data_out_0_79, E => ml_ms_output_edgedet, Q => ml_ms_sr11_data_out_1_80);
  ml_ms_sr11_data_out_reg_0 : EDFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_20, D => FE_PHN307_data_in, E => ml_ms_output_edgedet, Q => ml_ms_sr11_data_out_0_79);
  ml_ms_sr11_data_out_reg_3 : EDFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_20, D => FE_PHN279_ml_ms_data_sr_11bit_2, E => ml_ms_output_edgedet, Q => FE_PHN542_ml_ms_data_sr_11bit_3);
  ml_ms_sr11_data_out_reg_4 : EDFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_20, D => ml_ms_data_sr_11bit(3), E => ml_ms_output_edgedet, Q => FE_PHN90_ml_ms_data_sr_11bit_4);
  ml_ms_sr11_data_out_reg_5 : EDFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_20, D => ml_ms_data_sr_11bit(4), E => ml_ms_output_edgedet, Q => ml_ms_sr11_data_out_5_84);
  ml_ms_sr11_data_out_reg_7 : EDFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_20, D => ml_ms_data_sr_11bit(6), E => ml_ms_output_edgedet, Q => FE_PHN299_ml_ms_data_sr_11bit_7);
  ml_ms_sr11_data_out_reg_6 : EDFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_20, D => FE_PHN80_ml_ms_sr11_data_out_5_84, E => ml_ms_output_edgedet, Q => FE_PHN72_ml_ms_data_sr_11bit_6);
  ml_ms_sr11_data_out_reg_2 : EDFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_20, D => FE_PHN78_ml_ms_sr11_data_out_1_80, E => ml_ms_output_edgedet, Q => ml_ms_data_sr_11bit(2));
  ml_ms_flipflop4_Q_reg : DFXQD1BWP7T port map(CP => CTS_20, DA => ml_ms_mouse_y(0), DB => FE_PHN284_ml_mouseY_0, Q => ml_mouseY(0), SA => ml_ms_yflipfloprst);
  ml_ms_flipflop5_Q_reg : DFXQD1BWP7T port map(CP => CTS_20, DA => ml_ms_mouse_y(1), DB => FE_PHN79_ml_mouseY_1, Q => ml_mouseY(1), SA => ml_ms_yflipfloprst);
  ml_ms_flipflop6_Q_reg : DFXQD1BWP7T port map(CP => CTS_20, DA => ml_ms_mouse_y(2), DB => FE_PHN82_ml_mouseY_2, Q => ml_mouseY(2), SA => ml_ms_yflipfloprst);
  ml_ms_flipflop7_Q_reg : EDFQD1BWP7T port map(CP => CTS_20, D => ml_ms_btns(4), E => ml_ms_btnflipfloprst, Q => ml_buttons_mouse(4));
  ml_ms_flipflop8_Q_reg : DFXQD1BWP7T port map(CP => CTS_20, DA => ml_ms_btns(3), DB => FE_PHN320_ml_buttons_mouse_3, Q => ml_buttons_mouse(3), SA => ml_ms_btnflipfloprst);
  ml_ms_cnt_g71 : INVD1BWP7T port map(I => ml_ms_cntReset25M, ZN => ml_ms_cnt_n_23);
  ml_ms_cnt_count_reg_12 : DFKCNQD1BWP7T port map(CN => ml_ms_cnt_n_23, CP => CTS_20, D => FE_PHN368_ml_ms_cnt_n_22, Q => ml_ms_count25M(12));
  ml_ms_cnt_count_reg_11 : DFKCNQD1BWP7T port map(CN => ml_ms_cnt_n_23, CP => CTS_20, D => FE_PHN373_ml_ms_cnt_n_21, Q => ml_ms_count25M(11));
  ml_ms_cnt_g225 : MOAI22D0BWP7T port map(A1 => ml_ms_cnt_n_20, A2 => ml_ms_count25M(12), B1 => ml_ms_cnt_n_20, B2 => ml_ms_count25M(12), ZN => ml_ms_cnt_n_22);
  ml_ms_cnt_count_reg_10 : DFKCNQD1BWP7T port map(CN => ml_ms_cnt_n_23, CP => CTS_20, D => ml_ms_cnt_n_19, Q => ml_ms_count25M(10));
  ml_ms_cnt_g227 : MOAI22D0BWP7T port map(A1 => ml_ms_cnt_n_18, A2 => ml_ms_count25M(11), B1 => ml_ms_cnt_n_18, B2 => ml_ms_count25M(11), ZN => ml_ms_cnt_n_21);
  ml_ms_cnt_g228 : IND2D1BWP7T port map(A1 => ml_ms_cnt_n_18, B1 => ml_ms_count25M(11), ZN => ml_ms_cnt_n_20);
  ml_ms_cnt_count_reg_9 : DFKCNQD1BWP7T port map(CN => ml_ms_cnt_n_23, CP => CTS_20, D => ml_ms_cnt_n_17, Q => ml_ms_count25M(9));
  ml_ms_cnt_g230 : MOAI22D0BWP7T port map(A1 => ml_ms_cnt_n_16, A2 => ml_ms_count25M(10), B1 => ml_ms_cnt_n_16, B2 => ml_ms_count25M(10), ZN => FE_PHN363_ml_ms_cnt_n_19);
  ml_ms_cnt_g231 : IND2D1BWP7T port map(A1 => ml_ms_cnt_n_16, B1 => ml_ms_count25M(10), ZN => ml_ms_cnt_n_18);
  ml_ms_cnt_count_reg_8 : DFKCNQD1BWP7T port map(CN => ml_ms_cnt_n_23, CP => CTS_20, D => ml_ms_cnt_n_15, Q => FE_PHN452_ml_ms_count25M_8);
  ml_ms_cnt_g233 : MOAI22D0BWP7T port map(A1 => ml_ms_cnt_n_14, A2 => FE_PHN323_ml_ms_count25M_9, B1 => ml_ms_cnt_n_14, B2 => FE_PHN323_ml_ms_count25M_9, ZN => ml_ms_cnt_n_17);
  ml_ms_cnt_g234 : IND2D1BWP7T port map(A1 => ml_ms_cnt_n_14, B1 => FE_PHN323_ml_ms_count25M_9, ZN => ml_ms_cnt_n_16);
  ml_ms_cnt_count_reg_7 : DFKCNQD1BWP7T port map(CN => ml_ms_cnt_n_23, CP => CTS_20, D => ml_ms_cnt_n_13, Q => ml_ms_count25M(7));
  ml_ms_cnt_g236 : MOAI22D0BWP7T port map(A1 => ml_ms_cnt_n_12, A2 => ml_ms_count25M(8), B1 => ml_ms_cnt_n_12, B2 => ml_ms_count25M(8), ZN => ml_ms_cnt_n_15);
  ml_ms_cnt_g237 : IND2D1BWP7T port map(A1 => ml_ms_cnt_n_12, B1 => ml_ms_count25M(8), ZN => ml_ms_cnt_n_14);
  ml_ms_cnt_count_reg_6 : DFKCNQD1BWP7T port map(CN => ml_ms_cnt_n_11, CP => CTS_20, D => ml_ms_cnt_n_23, Q => ml_ms_count25M(6));
  ml_ms_cnt_g239 : MOAI22D0BWP7T port map(A1 => ml_ms_cnt_n_10, A2 => FE_PHN63_ml_ms_count25M_7, B1 => ml_ms_cnt_n_10, B2 => FE_PHN63_ml_ms_count25M_7, ZN => ml_ms_cnt_n_13);
  ml_ms_cnt_g240 : IND2D1BWP7T port map(A1 => ml_ms_cnt_n_10, B1 => FE_PHN63_ml_ms_count25M_7, ZN => ml_ms_cnt_n_12);
  ml_ms_cnt_count_reg_5 : DFKCNQD1BWP7T port map(CN => FE_PHN390_ml_ms_cnt_n_9, CP => CTS_20, D => ml_ms_cnt_n_23, Q => ml_ms_count25M(5));
  ml_ms_cnt_g242 : MOAI22D0BWP7T port map(A1 => ml_ms_cnt_n_8, A2 => FE_PHN318_ml_ms_count25M_6, B1 => ml_ms_cnt_n_8, B2 => FE_PHN318_ml_ms_count25M_6, ZN => ml_ms_cnt_n_11);
  ml_ms_cnt_g243 : IND2D1BWP7T port map(A1 => ml_ms_cnt_n_8, B1 => FE_PHN318_ml_ms_count25M_6, ZN => ml_ms_cnt_n_10);
  ml_ms_cnt_count_reg_4 : DFKCNQD1BWP7T port map(CN => FE_PHN386_ml_ms_cnt_n_7, CP => CTS_20, D => ml_ms_cnt_n_23, Q => ml_ms_count25M(4));
  ml_ms_cnt_g245 : MOAI22D0BWP7T port map(A1 => ml_ms_cnt_n_6, A2 => FE_PHN308_ml_ms_count25M_5, B1 => ml_ms_cnt_n_6, B2 => FE_PHN308_ml_ms_count25M_5, ZN => ml_ms_cnt_n_9);
  ml_ms_cnt_g246 : IND2D1BWP7T port map(A1 => ml_ms_cnt_n_6, B1 => FE_PHN308_ml_ms_count25M_5, ZN => ml_ms_cnt_n_8);
  ml_ms_cnt_count_reg_3 : DFKCNQD1BWP7T port map(CN => FE_PHN393_ml_ms_cnt_n_5, CP => CTS_20, D => ml_ms_cnt_n_23, Q => ml_ms_count25M(3));
  ml_ms_cnt_g248 : MOAI22D0BWP7T port map(A1 => ml_ms_cnt_n_4, A2 => ml_ms_count25M(4), B1 => ml_ms_cnt_n_4, B2 => ml_ms_count25M(4), ZN => ml_ms_cnt_n_7);
  ml_ms_cnt_g249 : IND2D1BWP7T port map(A1 => ml_ms_cnt_n_4, B1 => ml_ms_count25M(4), ZN => ml_ms_cnt_n_6);
  ml_ms_cnt_count_reg_2 : DFKCNQD1BWP7T port map(CN => FE_PHN383_ml_ms_cnt_n_3, CP => CTS_20, D => ml_ms_cnt_n_23, Q => ml_ms_count25M(2));
  ml_ms_cnt_g251 : MOAI22D0BWP7T port map(A1 => ml_ms_cnt_n_2, A2 => ml_ms_count25M(3), B1 => ml_ms_cnt_n_2, B2 => ml_ms_count25M(3), ZN => ml_ms_cnt_n_5);
  ml_ms_cnt_g252 : IND2D1BWP7T port map(A1 => ml_ms_cnt_n_2, B1 => ml_ms_count25M(3), ZN => ml_ms_cnt_n_4);
  ml_ms_cnt_count_reg_1 : EDFKCND1BWP7T port map(CN => ml_ms_cnt_n_23, CP => CTS_20, D => FE_PHN341_ml_ms_cnt_count_1, E => FE_PHN410_ml_ms_cnt_count_0, Q => UNCONNECTED0, QN => ml_ms_cnt_count(1));
  ml_ms_cnt_g254 : MOAI22D0BWP7T port map(A1 => ml_ms_cnt_n_1, A2 => ml_ms_count25M(2), B1 => ml_ms_cnt_n_1, B2 => ml_ms_count25M(2), ZN => ml_ms_cnt_n_3);
  ml_ms_cnt_g255 : IND2D1BWP7T port map(A1 => ml_ms_cnt_n_1, B1 => ml_ms_count25M(2), ZN => ml_ms_cnt_n_2);
  ml_ms_cnt_g257 : IND2D1BWP7T port map(A1 => FE_PHN341_ml_ms_cnt_count_1, B1 => ml_ms_cnt_count(0), ZN => ml_ms_cnt_n_1);
  ml_ms_cnt_count_reg_0 : DFKCND1BWP7T port map(CN => FE_PHN91_ml_ms_cnt_n_0, CP => CTS_20, D => ml_ms_cnt_n_23, Q => ml_ms_cnt_count(0), QN => ml_ms_cnt_n_0);
  ml_ms_flipflop9_Q_reg : EDFQD1BWP7T port map(CP => CTS_20, D => ml_ms_btns(2), E => ml_ms_btnflipfloprst, Q => ml_buttons_mouse(2));
  ml_ms_mx_g23 : ND2D5BWP7T port map(A1 => ml_ms_mx_n_0, A2 => ml_ms_mx_n_1, ZN => data_switch);
  ml_ms_mx_g24 : ND2D1BWP7T port map(A1 => FE_PHN446_ml_ms_mux_select, A2 => ml_ms_muxReg, ZN => ml_ms_mx_n_1);
  ml_ms_mx_g25 : IND2D1BWP7T port map(A1 => FE_PHN446_ml_ms_mux_select, B1 => FE_PHN526_ml_ms_muxFSM, ZN => ml_ms_mx_n_0);
  ml_ms_mx2_g23 : MUX2D1BWP7T port map(I0 => ml_ms_cntReset25M_main, I1 => ml_ms_cntReset25M_send, S => ml_ms_mux_select_main, Z => ml_ms_cntReset25M);
  ml_ms_cntD_g71 : INVD1BWP7T port map(I => FE_PHN68_ml_ms_count_debounce_reset, ZN => ml_ms_cntD_n_23);
  ml_ms_cntD_count_reg_12 : DFKCNQD1BWP7T port map(CN => ml_ms_cntD_n_23, CP => CTS_20, D => ml_ms_cntD_n_22, Q => ml_ms_count_debounce(12));
  ml_ms_cntD_count_reg_11 : DFKCNQD1BWP7T port map(CN => ml_ms_cntD_n_23, CP => CTS_20, D => ml_ms_cntD_n_21, Q => ml_ms_count_debounce(11));
  ml_ms_cntD_g225 : MOAI22D0BWP7T port map(A1 => ml_ms_cntD_n_20, A2 => FE_PHN666_ml_ms_count_debounce_12, B1 => ml_ms_cntD_n_20, B2 => FE_PHN663_ml_ms_count_debounce_12, ZN => ml_ms_cntD_n_22);
  ml_ms_cntD_count_reg_10 : DFKCNQD1BWP7T port map(CN => ml_ms_cntD_n_23, CP => CTS_20, D => FE_PHN397_ml_ms_cntD_n_19, Q => ml_ms_count_debounce(10));
  ml_ms_cntD_g227 : MOAI22D0BWP7T port map(A1 => ml_ms_cntD_n_18, A2 => FE_PHN123_ml_ms_count_debounce_11, B1 => ml_ms_cntD_n_18, B2 => FE_PHN123_ml_ms_count_debounce_11, ZN => ml_ms_cntD_n_21);
  ml_ms_cntD_g228 : IND2D1BWP7T port map(A1 => ml_ms_cntD_n_18, B1 => FE_PHN123_ml_ms_count_debounce_11, ZN => ml_ms_cntD_n_20);
  ml_ms_cntD_count_reg_9 : DFKCNQD1BWP7T port map(CN => ml_ms_cntD_n_23, CP => CTS_20, D => ml_ms_cntD_n_17, Q => ml_ms_count_debounce(9));
  ml_ms_cntD_g230 : MOAI22D0BWP7T port map(A1 => ml_ms_cntD_n_16, A2 => ml_ms_count_debounce(10), B1 => ml_ms_cntD_n_16, B2 => ml_ms_count_debounce(10), ZN => ml_ms_cntD_n_19);
  ml_ms_cntD_g231 : IND2D1BWP7T port map(A1 => ml_ms_cntD_n_16, B1 => FE_PHN617_ml_ms_count_debounce_10, ZN => ml_ms_cntD_n_18);
  ml_ms_cntD_count_reg_8 : DFKCNQD1BWP7T port map(CN => ml_ms_cntD_n_23, CP => CTS_20, D => ml_ms_cntD_n_15, Q => FE_PHN62_ml_ms_count_debounce_8);
  ml_ms_cntD_g233 : MOAI22D0BWP7T port map(A1 => ml_ms_cntD_n_14, A2 => FE_PHN61_ml_ms_count_debounce_9, B1 => ml_ms_cntD_n_14, B2 => FE_PHN61_ml_ms_count_debounce_9, ZN => ml_ms_cntD_n_17);
  ml_ms_cntD_g234 : IND2D1BWP7T port map(A1 => ml_ms_cntD_n_14, B1 => FE_PHN61_ml_ms_count_debounce_9, ZN => ml_ms_cntD_n_16);
  ml_ms_cntD_count_reg_7 : DFKCNQD1BWP7T port map(CN => ml_ms_cntD_n_23, CP => CTS_20, D => ml_ms_cntD_n_13, Q => ml_ms_count_debounce(7));
  ml_ms_cntD_g236 : MOAI22D0BWP7T port map(A1 => ml_ms_cntD_n_12, A2 => ml_ms_count_debounce(8), B1 => ml_ms_cntD_n_12, B2 => ml_ms_count_debounce(8), ZN => ml_ms_cntD_n_15);
  ml_ms_cntD_g237 : IND2D1BWP7T port map(A1 => ml_ms_cntD_n_12, B1 => ml_ms_count_debounce(8), ZN => ml_ms_cntD_n_14);
  ml_ms_cntD_count_reg_6 : DFKCNQD1BWP7T port map(CN => ml_ms_cntD_n_23, CP => CTS_20, D => ml_ms_cntD_n_11, Q => FE_PHN434_ml_ms_count_debounce_6);
  ml_ms_cntD_g239 : MOAI22D0BWP7T port map(A1 => ml_ms_cntD_n_10, A2 => FE_PHN473_ml_ms_count_debounce_7, B1 => ml_ms_cntD_n_10, B2 => FE_PHN473_ml_ms_count_debounce_7, ZN => ml_ms_cntD_n_13);
  ml_ms_cntD_g240 : IND2D1BWP7T port map(A1 => ml_ms_cntD_n_10, B1 => FE_PHN473_ml_ms_count_debounce_7, ZN => ml_ms_cntD_n_12);
  ml_ms_cntD_count_reg_5 : DFKCNQD1BWP7T port map(CN => ml_ms_cntD_n_23, CP => CTS_20, D => ml_ms_cntD_n_9, Q => ml_ms_count_debounce(5));
  ml_ms_cntD_g242 : MOAI22D0BWP7T port map(A1 => ml_ms_cntD_n_8, A2 => FE_PHN513_ml_ms_count_debounce_6, B1 => ml_ms_cntD_n_8, B2 => FE_PHN513_ml_ms_count_debounce_6, ZN => ml_ms_cntD_n_11);
  ml_ms_cntD_g243 : IND2D1BWP7T port map(A1 => ml_ms_cntD_n_8, B1 => FE_PHN513_ml_ms_count_debounce_6, ZN => ml_ms_cntD_n_10);
  ml_ms_cntD_count_reg_4 : DFKCNQD1BWP7T port map(CN => ml_ms_cntD_n_23, CP => CTS_20, D => ml_ms_cntD_n_7, Q => FE_PHN65_ml_ms_count_debounce_4);
  ml_ms_cntD_g245 : MOAI22D0BWP7T port map(A1 => ml_ms_cntD_n_6, A2 => FE_PHN69_ml_ms_count_debounce_5, B1 => ml_ms_cntD_n_6, B2 => FE_PHN69_ml_ms_count_debounce_5, ZN => ml_ms_cntD_n_9);
  ml_ms_cntD_g246 : IND2D1BWP7T port map(A1 => ml_ms_cntD_n_6, B1 => FE_PHN69_ml_ms_count_debounce_5, ZN => ml_ms_cntD_n_8);
  ml_ms_cntD_count_reg_3 : DFKCNQD1BWP7T port map(CN => ml_ms_cntD_n_23, CP => CTS_21, D => ml_ms_cntD_n_5, Q => FE_PHN64_ml_ms_count_debounce_3);
  ml_ms_cntD_g248 : MOAI22D0BWP7T port map(A1 => ml_ms_cntD_n_4, A2 => ml_ms_count_debounce(4), B1 => ml_ms_cntD_n_4, B2 => ml_ms_count_debounce(4), ZN => ml_ms_cntD_n_7);
  ml_ms_cntD_g249 : IND2D1BWP7T port map(A1 => ml_ms_cntD_n_4, B1 => ml_ms_count_debounce(4), ZN => ml_ms_cntD_n_6);
  ml_ms_cntD_count_reg_2 : DFKCNQD1BWP7T port map(CN => ml_ms_cntD_n_23, CP => CTS_21, D => ml_ms_cntD_n_3, Q => FE_PHN58_ml_ms_cntD_count_2);
  ml_ms_cntD_g251 : MOAI22D0BWP7T port map(A1 => ml_ms_cntD_n_2, A2 => ml_ms_count_debounce(3), B1 => ml_ms_cntD_n_2, B2 => ml_ms_count_debounce(3), ZN => ml_ms_cntD_n_5);
  ml_ms_cntD_g252 : IND2D1BWP7T port map(A1 => ml_ms_cntD_n_2, B1 => ml_ms_count_debounce(3), ZN => ml_ms_cntD_n_4);
  ml_ms_cntD_count_reg_1 : EDFKCND1BWP7T port map(CN => ml_ms_cntD_n_23, CP => CTS_20, D => ml_ms_cntD_count(1), E => FE_PHN60_ml_ms_cntD_count_0, Q => UNCONNECTED1, QN => FE_PHN313_ml_ms_cntD_count_1);
  ml_ms_cntD_g254 : MOAI22D0BWP7T port map(A1 => ml_ms_cntD_n_1, A2 => ml_ms_cntD_count(2), B1 => ml_ms_cntD_n_1, B2 => ml_ms_cntD_count(2), ZN => ml_ms_cntD_n_3);
  ml_ms_cntD_g255 : IND2D1BWP7T port map(A1 => ml_ms_cntD_n_1, B1 => ml_ms_cntD_count(2), ZN => ml_ms_cntD_n_2);
  ml_ms_cntD_g257 : IND2D1BWP7T port map(A1 => ml_ms_cntD_count(1), B1 => FE_PHN60_ml_ms_cntD_count_0, ZN => ml_ms_cntD_n_1);
  ml_ms_cntD_count_reg_0 : DFKCND1BWP7T port map(CN => FE_PHN89_ml_ms_cntD_n_0, CP => CTS_20, D => ml_ms_cntD_n_23, Q => ml_ms_cntD_count(0), QN => ml_ms_cntD_n_0);
  gl_const_gr_lg_mul_88_58_g474 : FA1D0BWP7T port map(A => gl_const_gr_lg_mul_88_58_n_7, B => gl_gr_lg_sig_countdown(10), CI => gl_const_gr_lg_mul_88_58_n_41, CO => gl_n_101, S => gl_n_100);
  gl_const_gr_lg_mul_88_58_g475 : FA1D0BWP7T port map(A => gl_const_gr_lg_mul_88_58_n_8, B => gl_const_gr_lg_mul_88_58_n_3, CI => gl_const_gr_lg_mul_88_58_n_39, CO => gl_const_gr_lg_mul_88_58_n_41, S => gl_n_99);
  gl_const_gr_lg_mul_88_58_g476 : FA1D0BWP7T port map(A => gl_const_gr_lg_mul_88_58_n_19, B => gl_const_gr_lg_mul_88_58_n_4, CI => gl_const_gr_lg_mul_88_58_n_37, CO => gl_const_gr_lg_mul_88_58_n_39, S => gl_n_98);
  gl_const_gr_lg_mul_88_58_g477 : FA1D0BWP7T port map(A => gl_const_gr_lg_mul_88_58_n_20, B => gl_const_gr_lg_mul_88_58_n_17, CI => gl_const_gr_lg_mul_88_58_n_35, CO => gl_const_gr_lg_mul_88_58_n_37, S => gl_n_97);
  gl_const_gr_lg_mul_88_58_g478 : FA1D0BWP7T port map(A => gl_const_gr_lg_mul_88_58_n_18, B => gl_const_gr_lg_mul_88_58_n_11, CI => gl_const_gr_lg_mul_88_58_n_33, CO => gl_const_gr_lg_mul_88_58_n_35, S => gl_n_96);
  gl_const_gr_lg_mul_88_58_g479 : FA1D0BWP7T port map(A => gl_const_gr_lg_mul_88_58_n_12, B => gl_const_gr_lg_mul_88_58_n_21, CI => gl_const_gr_lg_mul_88_58_n_31, CO => gl_const_gr_lg_mul_88_58_n_33, S => gl_n_95);
  gl_const_gr_lg_mul_88_58_g480 : FA1D0BWP7T port map(A => gl_const_gr_lg_mul_88_58_n_22, B => gl_const_gr_lg_mul_88_58_n_15, CI => gl_const_gr_lg_mul_88_58_n_29, CO => gl_const_gr_lg_mul_88_58_n_31, S => gl_n_94);
  gl_const_gr_lg_mul_88_58_g481 : FA1D0BWP7T port map(A => gl_const_gr_lg_mul_88_58_n_16, B => gl_const_gr_lg_mul_88_58_n_13, CI => gl_const_gr_lg_mul_88_58_n_27, CO => gl_const_gr_lg_mul_88_58_n_29, S => gl_n_93);
  gl_const_gr_lg_mul_88_58_g482 : FA1D0BWP7T port map(A => gl_const_gr_lg_mul_88_58_n_14, B => gl_const_gr_lg_mul_88_58_n_9, CI => gl_const_gr_lg_mul_88_58_n_25, CO => gl_const_gr_lg_mul_88_58_n_27, S => gl_n_92);
  gl_const_gr_lg_mul_88_58_g483 : FA1D0BWP7T port map(A => gl_const_gr_lg_mul_88_58_n_10, B => gl_const_gr_lg_mul_88_58_n_5, CI => gl_const_gr_lg_mul_88_58_n_23, CO => gl_const_gr_lg_mul_88_58_n_25, S => gl_n_91);
  gl_const_gr_lg_mul_88_58_g484 : FA1D0BWP7T port map(A => gl_const_gr_lg_mul_88_58_n_1, B => FE_PHN352_gl_gr_lg_sig_countdown_1, CI => gl_const_gr_lg_mul_88_58_n_6, CO => gl_const_gr_lg_mul_88_58_n_23, S => gl_n_90);
  gl_const_gr_lg_mul_88_58_g485 : FA1D0BWP7T port map(A => FE_PHN355_gl_gr_lg_sig_countdown_5, B => gl_gr_lg_sig_countdown(7), CI => gl_gr_lg_sig_countdown(4), CO => gl_const_gr_lg_mul_88_58_n_21, S => gl_const_gr_lg_mul_88_58_n_22);
  gl_const_gr_lg_mul_88_58_g486 : FA1D0BWP7T port map(A => gl_gr_lg_sig_countdown(8), B => gl_gr_lg_sig_countdown(10), CI => gl_gr_lg_sig_countdown(7), CO => gl_const_gr_lg_mul_88_58_n_19, S => gl_const_gr_lg_mul_88_58_n_20);
  gl_const_gr_lg_mul_88_58_g487 : FA1D0BWP7T port map(A => gl_gr_lg_sig_countdown(7), B => gl_gr_lg_sig_countdown(9), CI => gl_gr_lg_sig_countdown(6), CO => gl_const_gr_lg_mul_88_58_n_17, S => gl_const_gr_lg_mul_88_58_n_18);
  gl_const_gr_lg_mul_88_58_g488 : FA1D0BWP7T port map(A => gl_gr_lg_sig_countdown(3), B => gl_gr_lg_sig_countdown(6), CI => gl_gr_lg_sig_countdown(4), CO => gl_const_gr_lg_mul_88_58_n_15, S => gl_const_gr_lg_mul_88_58_n_16);
  gl_const_gr_lg_mul_88_58_g489 : FA1D0BWP7T port map(A => gl_gr_lg_sig_countdown(3), B => FE_PHN355_gl_gr_lg_sig_countdown_5, CI => FE_PHN354_gl_gr_lg_sig_countdown_2, CO => gl_const_gr_lg_mul_88_58_n_13, S => gl_const_gr_lg_mul_88_58_n_14);
  gl_const_gr_lg_mul_88_58_g490 : FA1D0BWP7T port map(A => gl_gr_lg_sig_countdown(6), B => gl_gr_lg_sig_countdown(8), CI => FE_PHN355_gl_gr_lg_sig_countdown_5, CO => gl_const_gr_lg_mul_88_58_n_11, S => gl_const_gr_lg_mul_88_58_n_12);
  gl_const_gr_lg_mul_88_58_g491 : FA1D0BWP7T port map(A => FE_PHN354_gl_gr_lg_sig_countdown_2, B => gl_gr_lg_sig_countdown(4), CI => FE_PHN352_gl_gr_lg_sig_countdown_1, CO => gl_const_gr_lg_mul_88_58_n_9, S => gl_const_gr_lg_mul_88_58_n_10);
  gl_const_gr_lg_mul_88_58_g492 : HA1D0BWP7T port map(A => gl_gr_lg_sig_countdown(9), B => gl_gr_lg_sig_countdown(10), CO => gl_const_gr_lg_mul_88_58_n_7, S => gl_const_gr_lg_mul_88_58_n_8);
  gl_const_gr_lg_mul_88_58_g493 : HA1D0BWP7T port map(A => gl_gr_lg_sig_countdown(3), B => FE_PHN353_gl_gr_lg_sig_countdown_0, CO => gl_const_gr_lg_mul_88_58_n_5, S => gl_const_gr_lg_mul_88_58_n_6);
  gl_const_gr_lg_mul_88_58_g494 : HA1D0BWP7T port map(A => gl_gr_lg_sig_countdown(9), B => gl_gr_lg_sig_countdown(8), CO => gl_const_gr_lg_mul_88_58_n_3, S => gl_const_gr_lg_mul_88_58_n_4);
  gl_const_gr_lg_mul_88_58_g495 : HA1D0BWP7T port map(A => gl_gr_lg_sig_countdown(2), B => FE_PHN353_gl_gr_lg_sig_countdown_0, CO => gl_const_gr_lg_mul_88_58_n_1, S => gl_n_89);
  gl_vga_buf_R1_Q_reg : EDFQD1BWP7T port map(CP => CTS_20, D => gl_Rint, E => FE_DBTN0_reset, Q => gl_vga_buf_Rint);
  gl_gr_lg_lh_l_edge_g12 : NR2XD0BWP7T port map(A1 => gl_gr_lg_lh_l_edge_n_0, A2 => gl_gr_lg_lh_l_edge_reg2, ZN => gl_gr_lg_lh_sig_edges);
  gl_gr_lg_lh_l_edge_reg2_reg : DFQD1BWP7T port map(CP => CTS_19, D => FE_PHN51_gl_gr_lg_lh_l_edge_reg1, Q => gl_gr_lg_lh_l_edge_reg2);
  gl_gr_lg_lh_l_edge_reg1_reg : DFD1BWP7T port map(CP => CTS_19, D => FE_PHN357_gl_sig_scale_h, Q => gl_gr_lg_lh_l_edge_reg1, QN => gl_gr_lg_lh_l_edge_n_0);
  gl_vga_buf_R2_Q_reg : EDFQD0BWP7T port map(CP => CTS_20, D => FE_PHN71_gl_vga_buf_Rint, E => FE_DBTN0_reset, Q => FE_OFN34_R);
  gl_gr_lg_lv_g307 : OAI32D1BWP7T port map(A1 => gl_gr_lg_local_y(2), A2 => gl_gr_lg_lv_n_5, A3 => gl_gr_lg_lv_n_8, B1 => FE_PHN407_gl_gr_lg_lv_n_3, B2 => gl_gr_lg_lv_n_13, ZN => gl_gr_lg_lv_n_15);
  gl_gr_lg_lv_g308 : OAI22D0BWP7T port map(A1 => gl_gr_lg_lv_n_13, A2 => gl_gr_lg_lv_n_4, B1 => gl_gr_lg_lv_n_8, B2 => gl_gr_lg_lv_n_11, ZN => gl_gr_lg_lv_n_14);
  gl_gr_lg_lv_count_v_reg_0 : DFXQD1BWP7T port map(CP => CTS_19, DA => gl_gr_lg_lv_n_10, DB => gl_gr_lg_lv_n_9, Q => FE_PHN348_gl_gr_lg_local_y_0, SA => FE_PHN465_gl_gr_lg_local_y_0);
  gl_gr_lg_lv_g311 : AOI21D0BWP7T port map(A1 => gl_gr_lg_lv_n_9, A2 => gl_gr_lg_lv_n_5, B => gl_gr_lg_lv_n_10, ZN => gl_gr_lg_lv_n_13);
  gl_gr_lg_lv_g312 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_lv_n_8, A2 => gl_gr_lg_lv_n_0, B1 => gl_gr_lg_lv_n_10, B2 => gl_gr_lg_local_y(1), ZN => gl_gr_lg_lv_n_12);
  gl_gr_lg_lv_g313 : OA32D1BWP7T port map(A1 => gl_gr_lg_local_y(3), A2 => gl_gr_lg_lv_n_3, A3 => gl_gr_lg_lv_n_5, B1 => gl_gr_lg_local_y(2), B2 => gl_gr_lg_lv_n_4, Z => gl_gr_lg_lv_n_11);
  gl_gr_lg_lv_g314 : NR2D1BWP7T port map(A1 => gl_gr_lg_lv_n_7, A2 => FE_PHN325_gl_gr_lg_lv_sig_edges, ZN => gl_gr_lg_lv_n_10);
  gl_gr_lg_lv_g315 : INVD0BWP7T port map(I => gl_gr_lg_lv_n_9, ZN => gl_gr_lg_lv_n_8);
  gl_gr_lg_lv_g316 : INR2XD0BWP7T port map(A1 => FE_PHN325_gl_gr_lg_lv_sig_edges, B1 => gl_gr_lg_lv_n_7, ZN => gl_gr_lg_lv_n_9);
  gl_gr_lg_lv_g317 : IND2D1BWP7T port map(A1 => FE_OFN35_reset, B1 => gl_gr_lg_lv_n_6, ZN => gl_gr_lg_lv_n_7);
  gl_gr_lg_lv_g318 : IND4D0BWP7T port map(A1 => gl_gr_lg_local_y(0), B1 => gl_gr_lg_local_y(3), B2 => gl_gr_lg_local_y(2), B3 => gl_gr_lg_local_y(1), ZN => gl_gr_lg_lv_n_6);
  gl_gr_lg_lv_g320 : ND2D1BWP7T port map(A1 => gl_gr_lg_local_y(1), A2 => gl_gr_lg_local_y(0), ZN => gl_gr_lg_lv_n_5);
  gl_gr_lg_lv_g2 : MUX2ND0BWP7T port map(I0 => gl_gr_lg_local_y(1), I1 => gl_gr_lg_lv_n_1, S => gl_gr_lg_local_y(0), ZN => gl_gr_lg_lv_n_0);
  gl_gr_lg_lv_count_v_reg_3 : DFD1BWP7T port map(CP => CTS_19, D => FE_PHN364_gl_gr_lg_lv_n_14, Q => gl_gr_lg_local_y(3), QN => gl_gr_lg_lv_n_4);
  gl_gr_lg_lv_count_v_reg_2 : DFD1BWP7T port map(CP => CTS_19, D => FE_PHN455_gl_gr_lg_lv_n_15, Q => gl_gr_lg_local_y(2), QN => gl_gr_lg_lv_n_3);
  gl_gr_lg_lv_count_v_reg_1 : DFD1BWP7T port map(CP => CTS_19, D => FE_PHN380_gl_gr_lg_lv_n_12, Q => gl_gr_lg_local_y(1), QN => gl_gr_lg_lv_n_1);
  gl_gr_lg_lv_l_edge_g12 : NR2XD0BWP7T port map(A1 => gl_gr_lg_lv_l_edge_n_0, A2 => gl_gr_lg_lv_l_edge_reg2, ZN => gl_gr_lg_lv_sig_edges);
  gl_gr_lg_lv_l_edge_reg2_reg : DFQD1BWP7T port map(CP => CTS_19, D => FE_PHN52_gl_gr_lg_lv_l_edge_reg1, Q => gl_gr_lg_lv_l_edge_reg2);
  gl_gr_lg_lv_l_edge_reg1_reg : DFD1BWP7T port map(CP => CTS_19, D => gl_sig_scale_v, Q => gl_gr_lg_lv_l_edge_reg1, QN => gl_gr_lg_lv_l_edge_n_0);
  ml_il_color1_g517 : INVD0BWP7T port map(I => sig_countlow, ZN => ml_il_color1_n_18);
  ml_il_color1_g591 : AO21D0BWP7T port map(A1 => sig_output_color(1), A2 => ml_il_color1_n_16, B => ml_il_color1_n_23, Z => sig_output_color(2));
  ml_il_color1_g592 : HA1D0BWP7T port map(A => ml_il_color1_state(1), B => ml_il_color1_state(2), CO => ml_il_color1_n_23, S => sig_output_color(1));
  ml_il_color1_g593 : OAI21D0BWP7T port map(A1 => ml_il_color1_n_17, A2 => ml_il_color1_state(1), B => ml_il_color1_n_24, ZN => sig_output_color(0));
  ml_il_color1_rescount_reg : DFKCNQD1BWP7T port map(CN => FE_PHN320_ml_buttons_mouse_3, CP => CTS_19, D => ml_il_color1_n_18, Q => sig_rescount);
  ml_il_color1_draw_reg : DFQD1BWP7T port map(CP => CTS_19, D => FE_PHN55_ml_buttons_mouse_4, Q => sig_draw);
  ml_il_color1_g596 : NR2D1BWP7T port map(A1 => ml_il_color1_state(2), A2 => ml_il_color1_state(0), ZN => ml_il_color1_n_17);
  ml_il_color1_g597 : ND2D1BWP7T port map(A1 => ml_il_color1_state(2), A2 => ml_il_color1_state(0), ZN => ml_il_color1_n_24);
  ml_il_color1_g797 : AO221D0BWP7T port map(A1 => ml_il_color1_n_9, A2 => ml_il_color1_n_3, B1 => ml_il_color1_n_23, B2 => FE_DBTN0_reset, C => ml_il_color1_n_11, Z => ml_il_color1_n_15);
  ml_il_color1_g799 : OAI211D1BWP7T port map(A1 => ml_il_color1_n_24, A2 => ml_il_color1_n_6, B => ml_il_color1_n_12, C => ml_il_color1_n_4, ZN => FE_PHN385_ml_il_color1_n_14);
  ml_il_color1_state_hs_reg_1 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_20, D => ml_il_color1_n_8, Q => FE_PHN406_ml_il_color1_state_hs_1);
  ml_il_color1_g801 : OAI22D0BWP7T port map(A1 => ml_il_color1_n_7, A2 => FE_OFN35_reset, B1 => ml_il_color1_n_6, B2 => FE_PHN59_ml_il_color1_n_1, ZN => ml_il_color1_n_13);
  ml_il_color1_g802 : IIND4D0BWP7T port map(A1 => sig_output_color(1), A2 => ml_il_color1_state(0), B1 => ml_il_color1_n_3, B2 => FE_DBTN0_reset, ZN => ml_il_color1_n_12);
  ml_il_color1_state_hs_reg_0 : DFKCNQD1BWP7T port map(CN => ml_il_color1_n_5, CP => CTS_20, D => ml_handshake_mouse_out, Q => ml_il_color1_state_hs(0));
  ml_il_color1_g804 : INVD1BWP7T port map(I => ml_il_color1_n_10, ZN => ml_il_color1_n_11);
  ml_il_color1_g805 : OAI22D0BWP7T port map(A1 => ml_il_color1_n_4, A2 => ml_il_color1_state(1), B1 => ml_il_color1_n_24, B2 => FE_OFN35_reset, ZN => ml_il_color1_n_9);
  ml_il_color1_g806 : IND3D1BWP7T port map(A1 => ml_il_color1_n_6, B1 => ml_il_color1_state(1), B2 => FE_PHN59_ml_il_color1_n_1, ZN => FE_PHN374_ml_il_color1_n_10);
  ml_il_color1_g807 : IAO21D0BWP7T port map(A1 => ml_handshake_mouse_out, A2 => FE_PHN87_ml_il_color1_state_hs_0, B => ml_il_color1_n_5, ZN => ml_il_color1_n_8);
  ml_il_color1_g808 : AOI32D1BWP7T port map(A1 => ml_il_color1_n_0, A2 => ml_il_color1_state(0), A3 => ml_il_color1_state(2), B1 => ml_il_color1_n_24, B2 => ml_il_color1_state(1), ZN => ml_il_color1_n_7);
  ml_il_color1_g809 : OR2D1BWP7T port map(A1 => ml_il_color1_n_3, A2 => FE_OFN35_reset, Z => ml_il_color1_n_6);
  ml_il_color1_g810 : NR3D0BWP7T port map(A1 => FE_PHN87_ml_il_color1_state_hs_0, A2 => ml_il_color1_state_hs(1), A3 => FE_OFN35_reset, ZN => ml_il_color1_n_5);
  ml_il_color1_g811 : ND3D0BWP7T port map(A1 => FE_PHN59_ml_il_color1_n_1, A2 => ml_il_color1_state(0), A3 => FE_DBTN0_reset, ZN => ml_il_color1_n_4);
  ml_il_color1_g812 : CKAN2D1BWP7T port map(A1 => FE_PHN87_ml_il_color1_state_hs_0, A2 => ml_buttons_mouse(2), Z => ml_il_color1_n_3);
  ml_il_color1_state_reg_0 : DFD1BWP7T port map(CP => CTS_20, D => ml_il_color1_n_14, Q => ml_il_color1_state(0), QN => ml_il_color1_n_16);
  ml_il_color1_state_reg_2 : DFKCND1BWP7T port map(CN => ml_il_color1_n_10, CP => CTS_20, D => FE_PHN378_ml_il_color1_n_13, Q => ml_il_color1_state(2), QN => ml_il_color1_n_1);
  ml_il_color1_state_reg_1 : DFD1BWP7T port map(CP => CTS_20, D => FE_PHN461_ml_il_color1_n_15, Q => ml_il_color1_state(1), QN => ml_il_color1_n_0);
  gl_vgd_g1598 : IND3D1BWP7T port map(A1 => gl_vgd_horizontal(8), B1 => gl_vgd_horizontal(9), B2 => gl_vgd_n_80, ZN => FE_PHN297_gl_Hint);
  gl_vgd_g1599 : AN2D0BWP7T port map(A1 => gl_sig_red, A2 => gl_vgd_n_79, Z => gl_Rint);
  gl_vgd_g1601 : AN2D0BWP7T port map(A1 => gl_sig_blue, A2 => gl_vgd_n_79, Z => gl_Bint);
  gl_vgd_g1602 : INR4D0BWP7T port map(A1 => gl_vgd_n_71, B1 => gl_vgd_horizontal(1), B2 => gl_vgd_horizontal(0), B3 => FE_PHN321_gl_vgd_n_77, ZN => gl_sig_scale_h);
  gl_vgd_g1603 : AOI31D0BWP7T port map(A1 => gl_vgd_n_74, A2 => gl_vgd_horizontal(5), A3 => gl_vgd_horizontal(7), B => gl_vgd_n_78, ZN => gl_vgd_n_80);
  gl_vgd_g1604 : OR4D1BWP7T port map(A1 => FE_PHN66_gl_vgd_vertical_9, A2 => gl_vgd_vertical(4), A3 => gl_vgd_n_69, A4 => gl_vgd_n_76, Z => gl_sig_v);
  gl_vgd_g1605 : IINR4D0BWP7T port map(A1 => gl_vgd_n_75, A2 => gl_vgd_n_69, B1 => gl_vgd_vertical(0), B2 => FE_PHN66_gl_vgd_vertical_9, ZN => FE_PHN358_gl_sig_scale_v);
  gl_vgd_g1607 : OAI31D0BWP7T port map(A1 => gl_vgd_horizontal(4), A2 => gl_vgd_horizontal(7), A3 => gl_vgd_n_72, B => gl_vgd_n_68, ZN => gl_vgd_n_78);
  gl_vgd_g1608 : INR3D0BWP7T port map(A1 => gl_vgd_n_69, B1 => FE_PHN66_gl_vgd_vertical_9, B2 => FE_PHN321_gl_vgd_n_77, ZN => gl_vgd_n_79);
  gl_vgd_g1609 : IND2D1BWP7T port map(A1 => gl_vgd_horizontal(9), B1 => gl_vgd_n_73, ZN => gl_vgd_n_77);
  gl_vgd_g1610 : IND3D1BWP7T port map(A1 => gl_vgd_n_67, B1 => gl_vgd_vertical(3), B2 => gl_vgd_n_70, ZN => gl_vgd_n_76);
  gl_vgd_g1611 : INR3D0BWP7T port map(A1 => gl_vgd_n_67, B1 => gl_vgd_vertical(4), B2 => gl_vgd_vertical(3), ZN => gl_vgd_n_75);
  gl_vgd_g1612 : IOA21D1BWP7T port map(A1 => gl_vgd_horizontal(1), A2 => gl_vgd_horizontal(0), B => gl_vgd_n_71, ZN => gl_vgd_n_74);
  gl_vgd_g1613 : ND4D0BWP7T port map(A1 => gl_vgd_horizontal(5), A2 => gl_vgd_horizontal(7), A3 => gl_vgd_horizontal(8), A4 => gl_vgd_horizontal(6), ZN => gl_vgd_n_73);
  gl_vgd_g1614 : AO211D0BWP7T port map(A1 => gl_vgd_horizontal(2), A2 => gl_vgd_horizontal(1), B => gl_vgd_horizontal(5), C => gl_vgd_horizontal(3), Z => gl_vgd_n_72);
  gl_vgd_g1615 : MUX2ND0BWP7T port map(I0 => gl_vgd_vertical(1), I1 => gl_vgd_vertical(2), S => gl_vgd_vertical(0), ZN => gl_vgd_n_70);
  gl_vgd_g1616 : NR3D0BWP7T port map(A1 => gl_vgd_horizontal(4), A2 => gl_vgd_horizontal(2), A3 => gl_vgd_horizontal(3), ZN => gl_vgd_n_71);
  gl_vgd_g1617 : MAOI22D0BWP7T port map(A1 => gl_vgd_horizontal(7), A2 => gl_vgd_horizontal(6), B1 => gl_vgd_horizontal(7), B2 => gl_vgd_horizontal(6), ZN => gl_vgd_n_68);
  gl_vgd_g1618 : ND4D0BWP7T port map(A1 => gl_vgd_vertical(5), A2 => gl_vgd_vertical(8), A3 => gl_vgd_vertical(7), A4 => gl_vgd_vertical(6), ZN => gl_vgd_n_69);
  gl_vgd_g1619 : NR2D1BWP7T port map(A1 => gl_vgd_vertical(1), A2 => gl_vgd_vertical(2), ZN => gl_vgd_n_67);
  gl_vgd_scale_horizontal_reg_8 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => FE_PHN524_gl_vgd_horizontal_counter_8, Q => gl_vgd_horizontal(8));
  gl_vgd_vertical_reg_4 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => FE_PHN324_gl_vgd_vertical_counter_4, Q => gl_vgd_vertical(4));
  gl_vgd_scale_horizontal_reg_3 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => gl_vgd_horizontal_counter(3), Q => gl_vgd_horizontal(3));
  gl_vgd_vertical_reg_3 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => gl_vgd_vertical_counter(3), Q => gl_vgd_vertical(3));
  gl_vgd_horizontal_reg_0 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => FE_PHN340_gl_vgd_horizontal_counter_0, Q => gl_vgd_horizontal(0));
  gl_vgd_vertical_reg_2 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => gl_vgd_vertical_counter(2), Q => gl_vgd_vertical(2));
  gl_vgd_vertical_reg_1 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => gl_vgd_vertical_counter(1), Q => gl_vgd_vertical(1));
  gl_vgd_horizontal_reg_6 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => gl_vgd_horizontal_counter(6), Q => gl_vgd_horizontal(6));
  gl_vgd_horizontal_reg_5 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => FE_PHN343_gl_vgd_horizontal_counter_5, Q => gl_vgd_horizontal(5));
  gl_vgd_scale_horizontal_reg_1 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => FE_PHN345_gl_vgd_horizontal_counter_1, Q => gl_vgd_horizontal(1));
  gl_vgd_scale_vertical_reg_8 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => FE_PHN57_gl_vgd_vertical_counter_8, Q => gl_vgd_vertical(8));
  gl_vgd_scale_vertical_reg_7 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => gl_vgd_vertical_counter(7), Q => gl_vgd_vertical(7));
  gl_vgd_scale_vertical_reg_6 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => gl_vgd_vertical_counter(6), Q => gl_vgd_vertical(6));
  gl_vgd_vertical_reg_5 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => FE_PHN326_gl_vgd_vertical_counter_5, Q => gl_vgd_vertical(5));
  gl_vgd_scale_horizontal_reg_4 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => gl_vgd_horizontal_counter(4), Q => gl_vgd_horizontal(4));
  gl_vgd_horizontal_reg_9 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => gl_vgd_horizontal_counter(9), Q => gl_vgd_horizontal(9));
  gl_vgd_scale_horizontal_reg_2 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => FE_PHN344_gl_vgd_horizontal_counter_2, Q => gl_vgd_horizontal(2));
  gl_vgd_vertical_reg_0 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => gl_vgd_vertical_counter(0), Q => gl_vgd_vertical(0));
  gl_vgd_scale_vertical_reg_9 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => gl_vgd_vertical_counter(9), Q => gl_vgd_vertical(9));
  gl_vgd_horizontal_reg_7 : DFKCNQD1BWP7T port map(CN => FE_DBTN0_reset, CP => CTS_19, D => FE_PHN529_gl_vgd_horizontal_counter_7, Q => gl_vgd_horizontal(7));
  gl_vgd_g2 : IND2D1BWP7T port map(A1 => gl_sig_green, B1 => gl_vgd_n_79, ZN => gl_Gint);
  gl_vgd_horizontal_counter_reg_0 : DFKCNQD1BWP7T port map(CN => gl_vgd_n_6, CP => CTS_19, D => gl_vgd_n_41, Q => gl_vgd_horizontal_counter(0));
  gl_vgd_horizontal_counter_reg_1 : DFKCNQD1BWP7T port map(CN => gl_vgd_n_19, CP => CTS_19, D => gl_vgd_n_41, Q => gl_vgd_horizontal_counter(1));
  gl_vgd_horizontal_counter_reg_2 : DFKCNQD1BWP7T port map(CN => gl_vgd_n_24, CP => CTS_19, D => gl_vgd_n_41, Q => gl_vgd_horizontal_counter(2));
  gl_vgd_horizontal_counter_reg_3 : DFKCNQD1BWP7T port map(CN => gl_vgd_n_29, CP => CTS_19, D => gl_vgd_n_41, Q => FE_PHN342_gl_vgd_horizontal_counter_3);
  gl_vgd_horizontal_counter_reg_4 : DFKCNQD1BWP7T port map(CN => gl_vgd_n_32, CP => CTS_19, D => gl_vgd_n_41, Q => FE_PHN346_gl_vgd_horizontal_counter_4);
  gl_vgd_horizontal_counter_reg_5 : DFKCNQD1BWP7T port map(CN => gl_vgd_n_37, CP => CTS_19, D => gl_vgd_n_41, Q => gl_vgd_horizontal_counter(5));
  gl_vgd_horizontal_counter_reg_6 : DFKCNQD1BWP7T port map(CN => gl_vgd_n_46, CP => CTS_19, D => gl_vgd_n_41, Q => FE_PHN543_gl_vgd_horizontal_counter_6);
  gl_vgd_horizontal_counter_reg_7 : DFKCNQD1BWP7T port map(CN => gl_vgd_n_56, CP => CTS_20, D => gl_vgd_n_41, Q => gl_vgd_horizontal_counter(7));
  gl_vgd_horizontal_counter_reg_8 : DFKCNQD1BWP7T port map(CN => gl_vgd_n_41, CP => CTS_20, D => gl_vgd_n_62, Q => gl_vgd_horizontal_counter(8));
  gl_vgd_horizontal_counter_reg_9 : DFKCNQD1BWP7T port map(CN => gl_vgd_n_41, CP => CTS_19, D => gl_vgd_n_65, Q => FE_PHN339_gl_vgd_horizontal_counter_9);
  gl_vgd_vertical_counter_reg_0 : DFXQD1BWP7T port map(CP => CTS_19, DA => gl_vgd_n_44, DB => gl_vgd_n_43, Q => FE_PHN336_gl_vgd_vertical_counter_0, SA => gl_vgd_vertical_counter(0));
  gl_vgd_vertical_counter_reg_1 : DFQD1BWP7T port map(CP => CTS_19, D => gl_vgd_n_51, Q => FE_PHN333_gl_vgd_vertical_counter_1);
  gl_vgd_vertical_counter_reg_2 : DFQD1BWP7T port map(CP => CTS_19, D => gl_vgd_n_52, Q => FE_PHN337_gl_vgd_vertical_counter_2);
  gl_vgd_vertical_counter_reg_3 : DFQD1BWP7T port map(CP => CTS_19, D => gl_vgd_n_49, Q => FE_PHN322_gl_vgd_vertical_counter_3);
  gl_vgd_vertical_counter_reg_4 : DFQD1BWP7T port map(CP => CTS_19, D => gl_vgd_n_54, Q => gl_vgd_vertical_counter(4));
  gl_vgd_vertical_counter_reg_5 : DFQD1BWP7T port map(CP => CTS_19, D => gl_vgd_n_53, Q => gl_vgd_vertical_counter(5));
  gl_vgd_vertical_counter_reg_6 : DFQD1BWP7T port map(CP => CTS_19, D => gl_vgd_n_50, Q => FE_PHN330_gl_vgd_vertical_counter_6);
  gl_vgd_vertical_counter_reg_7 : DFQD1BWP7T port map(CP => CTS_19, D => gl_vgd_n_57, Q => FE_PHN328_gl_vgd_vertical_counter_7);
  gl_vgd_vertical_counter_reg_9 : DFQD1BWP7T port map(CP => CTS_19, D => FE_PHN371_gl_vgd_n_64, Q => FE_PHN331_gl_vgd_vertical_counter_9);
  gl_vgd_g1735 : MOAI22D0BWP7T port map(A1 => gl_vgd_n_63, A2 => gl_vgd_n_14, B1 => gl_vgd_n_63, B2 => gl_vgd_n_14, ZN => gl_vgd_n_65);
  gl_vgd_g1738 : AO22D0BWP7T port map(A1 => gl_vgd_n_58, A2 => gl_vgd_vertical_counter(9), B1 => gl_vgd_n_60, B2 => gl_vgd_n_43, Z => gl_vgd_n_64);
  gl_vgd_g1739 : HA1D0BWP7T port map(A => gl_vgd_n_11, B => gl_vgd_n_55, CO => gl_vgd_n_63, S => gl_vgd_n_62);
  gl_vgd_g1740 : AO21D0BWP7T port map(A1 => gl_vgd_n_58, A2 => FE_PHN57_gl_vgd_vertical_counter_8, B => gl_vgd_n_59, Z => gl_vgd_n_61);
  gl_vgd_g1742 : OAI31D0BWP7T port map(A1 => gl_vgd_vertical_counter(9), A2 => gl_vgd_n_2, A3 => gl_vgd_n_47, B => gl_vgd_n_15, ZN => gl_vgd_n_60);
  gl_vgd_g1744 : NR3D0BWP7T port map(A1 => gl_vgd_n_42, A2 => gl_vgd_n_47, A3 => FE_PHN57_gl_vgd_vertical_counter_8, ZN => gl_vgd_n_59);
  gl_vgd_g1745 : MOAI22D0BWP7T port map(A1 => gl_vgd_n_42, A2 => gl_vgd_n_48, B1 => gl_vgd_n_44, B2 => gl_vgd_vertical_counter(7), ZN => gl_vgd_n_57);
  gl_vgd_g1746 : AO21D0BWP7T port map(A1 => gl_vgd_n_43, A2 => gl_vgd_n_47, B => gl_vgd_n_44, Z => gl_vgd_n_58);
  gl_vgd_g1747 : HA1D0BWP7T port map(A => gl_vgd_n_13, B => gl_vgd_n_45, CO => gl_vgd_n_55, S => gl_vgd_n_56);
  gl_vgd_g1755 : MOAI22D0BWP7T port map(A1 => gl_vgd_n_42, A2 => gl_vgd_n_30, B1 => gl_vgd_n_44, B2 => FE_PHN324_gl_vgd_vertical_counter_4, ZN => gl_vgd_n_54);
  gl_vgd_g1756 : MOAI22D0BWP7T port map(A1 => gl_vgd_n_42, A2 => gl_vgd_n_34, B1 => gl_vgd_n_44, B2 => FE_PHN326_gl_vgd_vertical_counter_5, ZN => gl_vgd_n_53);
  gl_vgd_g1758 : MOAI22D0BWP7T port map(A1 => gl_vgd_n_42, A2 => gl_vgd_n_20, B1 => gl_vgd_n_44, B2 => gl_vgd_vertical_counter(2), ZN => gl_vgd_n_52);
  gl_vgd_g1759 : MOAI22D0BWP7T port map(A1 => gl_vgd_n_42, A2 => gl_vgd_n_0, B1 => gl_vgd_n_44, B2 => gl_vgd_vertical_counter(1), ZN => gl_vgd_n_51);
  gl_vgd_g1760 : MOAI22D0BWP7T port map(A1 => gl_vgd_n_42, A2 => gl_vgd_n_39, B1 => gl_vgd_n_44, B2 => gl_vgd_vertical_counter(6), ZN => gl_vgd_n_50);
  gl_vgd_g1761 : MOAI22D0BWP7T port map(A1 => gl_vgd_n_42, A2 => gl_vgd_n_25, B1 => gl_vgd_n_44, B2 => gl_vgd_vertical_counter(3), ZN => gl_vgd_n_49);
  gl_vgd_g1765 : MAOI22D0BWP7T port map(A1 => gl_vgd_n_38, A2 => gl_vgd_vertical_counter(7), B1 => gl_vgd_n_38, B2 => gl_vgd_vertical_counter(7), ZN => gl_vgd_n_48);
  gl_vgd_g1769 : HA1D0BWP7T port map(A => gl_vgd_n_12, B => gl_vgd_n_36, CO => gl_vgd_n_45, S => gl_vgd_n_46);
  gl_vgd_g1770 : IND2D1BWP7T port map(A1 => gl_vgd_n_38, B1 => gl_vgd_vertical_counter(7), ZN => gl_vgd_n_47);
  gl_vgd_g1771 : INVD1BWP7T port map(I => gl_vgd_n_43, ZN => gl_vgd_n_42);
  gl_vgd_g1772 : NR2D1BWP7T port map(A1 => gl_vgd_n_40, A2 => FE_OFN35_reset, ZN => gl_vgd_n_44);
  gl_vgd_g1773 : NR2XD0BWP7T port map(A1 => gl_vgd_n_41, A2 => gl_vgd_n_26, ZN => gl_vgd_n_43);
  gl_vgd_g1774 : INVD1BWP7T port map(I => gl_vgd_n_41, ZN => gl_vgd_n_40);
  gl_vgd_g1775 : IND3D1BWP7T port map(A1 => gl_vgd_n_13, B1 => gl_vgd_n_11, B2 => gl_vgd_n_35, ZN => gl_vgd_n_41);
  gl_vgd_g1776 : MAOI22D0BWP7T port map(A1 => gl_vgd_n_31, A2 => gl_vgd_vertical_counter(6), B1 => gl_vgd_n_31, B2 => gl_vgd_vertical_counter(6), ZN => gl_vgd_n_39);
  gl_vgd_g1777 : HA1D0BWP7T port map(A => gl_vgd_n_8, B => gl_vgd_n_33, CO => gl_vgd_n_36, S => gl_vgd_n_37);
  gl_vgd_g1778 : IND2D1BWP7T port map(A1 => gl_vgd_n_31, B1 => gl_vgd_vertical_counter(6), ZN => gl_vgd_n_38);
  gl_vgd_g1779 : INR4D0BWP7T port map(A1 => gl_vgd_n_33, B1 => gl_vgd_n_14, B2 => gl_vgd_n_8, B3 => gl_vgd_n_12, ZN => gl_vgd_n_35);
  gl_vgd_g1780 : MAOI22D0BWP7T port map(A1 => gl_vgd_n_27, A2 => FE_PHN326_gl_vgd_vertical_counter_5, B1 => gl_vgd_n_27, B2 => FE_PHN326_gl_vgd_vertical_counter_5, ZN => gl_vgd_n_34);
  gl_vgd_g1781 : HA1D0BWP7T port map(A => gl_vgd_n_10, B => gl_vgd_n_28, CO => gl_vgd_n_33, S => gl_vgd_n_32);
  gl_vgd_g1782 : IND2D1BWP7T port map(A1 => gl_vgd_n_27, B1 => FE_PHN326_gl_vgd_vertical_counter_5, ZN => gl_vgd_n_31);
  gl_vgd_g1783 : MAOI22D0BWP7T port map(A1 => gl_vgd_n_22, A2 => FE_PHN324_gl_vgd_vertical_counter_4, B1 => gl_vgd_n_22, B2 => FE_PHN324_gl_vgd_vertical_counter_4, ZN => gl_vgd_n_30);
  gl_vgd_g1784 : HA1D0BWP7T port map(A => gl_vgd_n_4, B => gl_vgd_n_23, CO => gl_vgd_n_28, S => gl_vgd_n_29);
  gl_vgd_g1785 : IND2D1BWP7T port map(A1 => gl_vgd_n_22, B1 => FE_PHN324_gl_vgd_vertical_counter_4, ZN => gl_vgd_n_27);
  gl_vgd_g1786 : NR4D0BWP7T port map(A1 => gl_vgd_n_21, A2 => gl_vgd_vertical_counter(7), A3 => gl_vgd_vertical_counter(6), A4 => FE_PHN326_gl_vgd_vertical_counter_5, ZN => gl_vgd_n_26);
  gl_vgd_g1787 : MAOI22D0BWP7T port map(A1 => gl_vgd_n_17, A2 => gl_vgd_vertical_counter(3), B1 => gl_vgd_n_17, B2 => gl_vgd_vertical_counter(3), ZN => gl_vgd_n_25);
  gl_vgd_g1788 : HA1D0BWP7T port map(A => gl_vgd_n_3, B => gl_vgd_n_18, CO => gl_vgd_n_23, S => gl_vgd_n_24);
  gl_vgd_g1789 : IND2D1BWP7T port map(A1 => gl_vgd_n_17, B1 => gl_vgd_vertical_counter(3), ZN => gl_vgd_n_22);
  gl_vgd_g1790 : IND4D0BWP7T port map(A1 => FE_PHN324_gl_vgd_vertical_counter_4, B1 => gl_vgd_vertical_counter(2), B2 => gl_vgd_vertical_counter(3), B3 => gl_vgd_n_16, ZN => gl_vgd_n_21);
  gl_vgd_g1791 : MAOI22D0BWP7T port map(A1 => gl_vgd_n_9, A2 => gl_vgd_vertical_counter(2), B1 => gl_vgd_n_9, B2 => gl_vgd_vertical_counter(2), ZN => gl_vgd_n_20);
  gl_vgd_g1792 : HA1D0BWP7T port map(A => gl_vgd_n_7, B => gl_vgd_n_5, CO => gl_vgd_n_18, S => gl_vgd_n_19);
  gl_vgd_g1793 : IND2D1BWP7T port map(A1 => gl_vgd_n_9, B1 => gl_vgd_vertical_counter(2), ZN => gl_vgd_n_17);
  gl_vgd_g1794 : NR3D0BWP7T port map(A1 => gl_vgd_n_15, A2 => gl_vgd_vertical_counter(1), A3 => gl_vgd_vertical_counter(0), ZN => gl_vgd_n_16);
  gl_vgd_g1796 : ND2D1BWP7T port map(A1 => gl_vgd_n_2, A2 => gl_vgd_vertical_counter(9), ZN => gl_vgd_n_15);
  gl_vgd_g1797 : ND2D1BWP7T port map(A1 => gl_vgd_horizontal_counter(9), A2 => FE_DBTN0_reset, ZN => gl_vgd_n_14);
  gl_vgd_g1798 : INR2XD0BWP7T port map(A1 => gl_vgd_horizontal_counter(4), B1 => FE_OFN35_reset, ZN => gl_vgd_n_10);
  gl_vgd_g1799 : INR2D1BWP7T port map(A1 => FE_PHN529_gl_vgd_horizontal_counter_7, B1 => FE_OFN35_reset, ZN => gl_vgd_n_13);
  gl_vgd_g1800 : INR2D1BWP7T port map(A1 => gl_vgd_horizontal_counter(6), B1 => FE_OFN35_reset, ZN => gl_vgd_n_12);
  gl_vgd_g1801 : INR2D1BWP7T port map(A1 => FE_PHN524_gl_vgd_horizontal_counter_8, B1 => FE_OFN35_reset, ZN => gl_vgd_n_11);
  gl_vgd_g1802 : INVD0BWP7T port map(I => gl_vgd_n_6, ZN => gl_vgd_n_7);
  gl_vgd_g1803 : CKAN2D1BWP7T port map(A1 => FE_PHN345_gl_vgd_horizontal_counter_1, A2 => FE_DBTN0_reset, Z => gl_vgd_n_5);
  gl_vgd_g1804 : ND2D1BWP7T port map(A1 => gl_vgd_vertical_counter(1), A2 => gl_vgd_vertical_counter(0), ZN => gl_vgd_n_9);
  gl_vgd_g1805 : CKAN2D1BWP7T port map(A1 => gl_vgd_horizontal_counter(3), A2 => FE_DBTN0_reset, Z => gl_vgd_n_4);
  gl_vgd_g1806 : CKAN2D1BWP7T port map(A1 => FE_PHN344_gl_vgd_horizontal_counter_2, A2 => FE_DBTN0_reset, Z => gl_vgd_n_3);
  gl_vgd_g1807 : AN2D1BWP7T port map(A1 => FE_PHN343_gl_vgd_horizontal_counter_5, A2 => FE_DBTN0_reset, Z => gl_vgd_n_8);
  gl_vgd_g1808 : ND2D1BWP7T port map(A1 => FE_PHN340_gl_vgd_horizontal_counter_0, A2 => FE_DBTN0_reset, ZN => gl_vgd_n_6);
  gl_vgd_g1641 : XNR2D1BWP7T port map(A1 => gl_vgd_vertical_counter(1), A2 => gl_vgd_vertical_counter(0), ZN => gl_vgd_n_0);
  gl_vgd_vertical_counter_reg_8 : DFD1BWP7T port map(CP => CTS_19, D => gl_vgd_n_61, Q => gl_vgd_vertical_counter(8), QN => gl_vgd_n_2);
  gl_gr_lg_div_88_62_g3670 : OAI22D0BWP7T port map(A1 => gl_n_84, A2 => gl_gr_lg_div_88_62_n_136, B1 => gl_gr_lg_div_88_62_n_137, B2 => gl_gr_lg_div_88_62_n_135, ZN => gl_n_85);
  gl_gr_lg_div_88_62_g3671 : OAI21D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_134, A2 => gl_gr_lg_div_88_62_n_131, B => gl_gr_lg_div_88_62_n_135, ZN => gl_n_84);
  gl_gr_lg_div_88_62_g3672 : NR4D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_128, A2 => gl_gr_lg_div_88_62_n_130, A3 => FE_PHN352_gl_gr_lg_sig_countdown_1, A4 => FE_PHN353_gl_gr_lg_sig_countdown_0, ZN => gl_gr_lg_div_88_62_n_137);
  gl_gr_lg_div_88_62_g3673 : AOI211XD0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_133, A2 => gl_gr_lg_div_88_62_n_130, B => gl_gr_lg_div_88_62_n_127, C => gl_gr_lg_div_88_62_n_125, ZN => gl_gr_lg_div_88_62_n_136);
  gl_gr_lg_div_88_62_g3674 : AOI21D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_132, A2 => gl_gr_lg_div_88_62_n_105, B => gl_gr_lg_div_88_62_n_129, ZN => gl_gr_lg_div_88_62_n_135);
  gl_gr_lg_div_88_62_g3675 : AOI21D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_128, A2 => FE_PHN352_gl_gr_lg_sig_countdown_1, B => gl_gr_lg_div_88_62_n_130, ZN => gl_gr_lg_div_88_62_n_134);
  gl_gr_lg_div_88_62_g3676 : AO21D0BWP7T port map(A1 => FE_PHN353_gl_gr_lg_sig_countdown_0, A2 => FE_PHN352_gl_gr_lg_sig_countdown_1, B => gl_gr_lg_div_88_62_n_128, Z => gl_gr_lg_div_88_62_n_133);
  gl_gr_lg_div_88_62_g3677 : OAI221D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_119, A2 => gl_gr_lg_div_88_62_n_114, B1 => gl_gr_lg_div_88_62_n_110, B2 => gl_gr_lg_div_88_62_n_121, C => gl_gr_lg_div_88_62_n_116, ZN => gl_gr_lg_div_88_62_n_132);
  gl_gr_lg_div_88_62_g3678 : NR2D1BWP7T port map(A1 => gl_gr_lg_div_88_62_n_127, A2 => gl_gr_lg_div_88_62_n_125, ZN => gl_gr_lg_div_88_62_n_131);
  gl_gr_lg_div_88_62_g3679 : OAI221D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_121, A2 => gl_n_90, B1 => gl_gr_lg_div_88_62_n_17, B2 => gl_gr_lg_div_88_62_n_119, C => gl_gr_lg_div_88_62_n_126, ZN => gl_gr_lg_div_88_62_n_130);
  gl_gr_lg_div_88_62_g3680 : OAI32D1BWP7T port map(A1 => gl_gr_lg_div_88_62_n_105, A2 => gl_gr_lg_div_88_62_n_109, A3 => gl_gr_lg_div_88_62_n_123, B1 => gl_gr_lg_div_88_62_n_117, B2 => gl_gr_lg_div_88_62_n_121, ZN => gl_gr_lg_div_88_62_n_129);
  gl_gr_lg_div_88_62_g3681 : MOAI22D0BWP7T port map(A1 => gl_n_86, A2 => gl_gr_lg_div_88_62_n_5, B1 => gl_n_86, B2 => gl_gr_lg_div_88_62_n_5, ZN => gl_gr_lg_div_88_62_n_128);
  gl_gr_lg_div_88_62_g3682 : OAI22D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_119, A2 => gl_gr_lg_div_88_62_n_113, B1 => gl_gr_lg_div_88_62_n_123, B2 => gl_gr_lg_div_88_62_n_118, ZN => gl_gr_lg_div_88_62_n_127);
  gl_gr_lg_div_88_62_g3683 : AOI22D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_115, A2 => gl_n_90, B1 => gl_gr_lg_div_88_62_n_122, B2 => gl_gr_lg_div_88_62_n_17, ZN => gl_gr_lg_div_88_62_n_126);
  gl_gr_lg_div_88_62_g3684 : OAI22D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_116, A2 => gl_gr_lg_div_88_62_n_102, B1 => gl_gr_lg_div_88_62_n_121, B2 => gl_gr_lg_div_88_62_n_111, ZN => gl_gr_lg_div_88_62_n_125);
  gl_gr_lg_div_88_62_g3685 : AN2D1BWP7T port map(A1 => gl_gr_lg_div_88_62_n_121, A2 => gl_gr_lg_div_88_62_n_116, Z => gl_n_86);
  gl_gr_lg_div_88_62_g3686 : INVD0BWP7T port map(I => gl_gr_lg_div_88_62_n_122, ZN => gl_gr_lg_div_88_62_n_123);
  gl_gr_lg_div_88_62_g3687 : NR2XD0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_115, A2 => gl_n_87, ZN => gl_gr_lg_div_88_62_n_122);
  gl_gr_lg_div_88_62_g3688 : ND2D1BWP7T port map(A1 => gl_n_87, A2 => gl_gr_lg_div_88_62_n_119, ZN => gl_gr_lg_div_88_62_n_121);
  gl_gr_lg_div_88_62_g3689 : IOA21D1BWP7T port map(A1 => gl_gr_lg_div_88_62_n_117, A2 => gl_gr_lg_div_88_62_n_107, B => gl_gr_lg_div_88_62_n_112, ZN => gl_n_87);
  gl_gr_lg_div_88_62_g3690 : AO21D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_114, A2 => gl_gr_lg_div_88_62_n_104, B => gl_gr_lg_div_88_62_n_112, Z => gl_gr_lg_div_88_62_n_119);
  gl_gr_lg_div_88_62_g3691 : IAO21D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_110, A2 => gl_gr_lg_div_88_62_n_5, B => gl_gr_lg_div_88_62_n_109, ZN => gl_gr_lg_div_88_62_n_118);
  gl_gr_lg_div_88_62_g3692 : ND2D1BWP7T port map(A1 => gl_gr_lg_div_88_62_n_110, A2 => gl_gr_lg_div_88_62_n_104, ZN => gl_gr_lg_div_88_62_n_117);
  gl_gr_lg_div_88_62_g3693 : INVD0BWP7T port map(I => gl_gr_lg_div_88_62_n_116, ZN => gl_gr_lg_div_88_62_n_115);
  gl_gr_lg_div_88_62_g3694 : OAI211D1BWP7T port map(A1 => gl_gr_lg_div_88_62_n_104, A2 => gl_gr_lg_div_88_62_n_109, B => gl_gr_lg_div_88_62_n_112, C => gl_gr_lg_div_88_62_n_108, ZN => gl_gr_lg_div_88_62_n_116);
  gl_gr_lg_div_88_62_g3695 : HA1D0BWP7T port map(A => gl_gr_lg_div_88_62_n_13, B => gl_gr_lg_div_88_62_n_102, CO => gl_gr_lg_div_88_62_n_114, S => gl_gr_lg_div_88_62_n_113);
  gl_gr_lg_div_88_62_g3696 : AOI21D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_106, A2 => gl_gr_lg_div_88_62_n_81, B => gl_gr_lg_div_88_62_n_103, ZN => gl_gr_lg_div_88_62_n_112);
  gl_gr_lg_div_88_62_g3697 : MAOI22D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_102, A2 => gl_n_90, B1 => gl_gr_lg_div_88_62_n_102, B2 => gl_n_90, ZN => gl_gr_lg_div_88_62_n_111);
  gl_gr_lg_div_88_62_g3698 : IND2D1BWP7T port map(A1 => gl_gr_lg_div_88_62_n_102, B1 => gl_n_90, ZN => gl_gr_lg_div_88_62_n_110);
  gl_gr_lg_div_88_62_g3699 : AOI21D0BWP7T port map(A1 => gl_n_90, A2 => gl_n_89, B => gl_gr_lg_div_88_62_n_101, ZN => gl_gr_lg_div_88_62_n_109);
  gl_gr_lg_div_88_62_g3700 : INVD0BWP7T port map(I => gl_gr_lg_div_88_62_n_107, ZN => gl_gr_lg_div_88_62_n_108);
  gl_gr_lg_div_88_62_g3701 : OAI221D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_95, A2 => gl_gr_lg_div_88_62_n_85, B1 => gl_gr_lg_div_88_62_n_77, B2 => gl_gr_lg_div_88_62_n_90, C => gl_gr_lg_div_88_62_n_100, ZN => gl_gr_lg_div_88_62_n_107);
  gl_gr_lg_div_88_62_g3702 : OAI221D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_95, A2 => gl_gr_lg_div_88_62_n_84, B1 => gl_gr_lg_div_88_62_n_88, B2 => gl_gr_lg_div_88_62_n_93, C => gl_gr_lg_div_88_62_n_90, ZN => gl_gr_lg_div_88_62_n_106);
  gl_gr_lg_div_88_62_g3703 : INVD1BWP7T port map(I => gl_gr_lg_div_88_62_n_105, ZN => gl_gr_lg_div_88_62_n_104);
  gl_gr_lg_div_88_62_g3704 : OAI221D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_95, A2 => gl_n_92, B1 => gl_gr_lg_div_88_62_n_16, B2 => gl_gr_lg_div_88_62_n_93, C => gl_gr_lg_div_88_62_n_99, ZN => gl_gr_lg_div_88_62_n_105);
  gl_gr_lg_div_88_62_g3705 : OAI32D1BWP7T port map(A1 => gl_gr_lg_div_88_62_n_81, A2 => gl_gr_lg_div_88_62_n_83, A3 => gl_gr_lg_div_88_62_n_97, B1 => gl_gr_lg_div_88_62_n_91, B2 => gl_gr_lg_div_88_62_n_95, ZN => gl_gr_lg_div_88_62_n_103);
  gl_gr_lg_div_88_62_g3706 : INVD0BWP7T port map(I => gl_gr_lg_div_88_62_n_102, ZN => gl_gr_lg_div_88_62_n_101);
  gl_gr_lg_div_88_62_g3707 : MAOI22D0BWP7T port map(A1 => gl_n_103, A2 => gl_gr_lg_div_88_62_n_4, B1 => gl_n_103, B2 => gl_gr_lg_div_88_62_n_4, ZN => gl_gr_lg_div_88_62_n_102);
  gl_gr_lg_div_88_62_g3708 : OA22D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_97, A2 => gl_gr_lg_div_88_62_n_92, B1 => gl_gr_lg_div_88_62_n_87, B2 => gl_gr_lg_div_88_62_n_93, Z => gl_gr_lg_div_88_62_n_100);
  gl_gr_lg_div_88_62_g3709 : AOI22D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_96, A2 => gl_gr_lg_div_88_62_n_16, B1 => gl_gr_lg_div_88_62_n_89, B2 => gl_n_92, ZN => gl_gr_lg_div_88_62_n_99);
  gl_gr_lg_div_88_62_g3710 : CKAN2D1BWP7T port map(A1 => gl_gr_lg_div_88_62_n_95, A2 => gl_gr_lg_div_88_62_n_90, Z => gl_n_103);
  gl_gr_lg_div_88_62_g3711 : INVD0BWP7T port map(I => gl_gr_lg_div_88_62_n_96, ZN => gl_gr_lg_div_88_62_n_97);
  gl_gr_lg_div_88_62_g3712 : NR2D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_89, A2 => gl_n_102, ZN => gl_gr_lg_div_88_62_n_96);
  gl_gr_lg_div_88_62_g3713 : ND2D1BWP7T port map(A1 => gl_n_102, A2 => gl_gr_lg_div_88_62_n_93, ZN => gl_gr_lg_div_88_62_n_95);
  gl_gr_lg_div_88_62_g3714 : IOA21D1BWP7T port map(A1 => gl_gr_lg_div_88_62_n_91, A2 => gl_gr_lg_div_88_62_n_79, B => gl_gr_lg_div_88_62_n_86, ZN => gl_n_102);
  gl_gr_lg_div_88_62_g3715 : AO21D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_88, A2 => gl_gr_lg_div_88_62_n_82, B => gl_gr_lg_div_88_62_n_86, Z => gl_gr_lg_div_88_62_n_93);
  gl_gr_lg_div_88_62_g3716 : IAO21D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_84, A2 => gl_gr_lg_div_88_62_n_4, B => gl_gr_lg_div_88_62_n_83, ZN => gl_gr_lg_div_88_62_n_92);
  gl_gr_lg_div_88_62_g3717 : ND2D1BWP7T port map(A1 => gl_gr_lg_div_88_62_n_84, A2 => gl_gr_lg_div_88_62_n_82, ZN => gl_gr_lg_div_88_62_n_91);
  gl_gr_lg_div_88_62_g3718 : INVD0BWP7T port map(I => gl_gr_lg_div_88_62_n_90, ZN => gl_gr_lg_div_88_62_n_89);
  gl_gr_lg_div_88_62_g3719 : OAI211D1BWP7T port map(A1 => gl_gr_lg_div_88_62_n_82, A2 => gl_gr_lg_div_88_62_n_83, B => gl_gr_lg_div_88_62_n_86, C => gl_gr_lg_div_88_62_n_78, ZN => gl_gr_lg_div_88_62_n_90);
  gl_gr_lg_div_88_62_g3720 : HA1D0BWP7T port map(A => gl_gr_lg_div_88_62_n_12, B => gl_gr_lg_div_88_62_n_77, CO => gl_gr_lg_div_88_62_n_88, S => gl_gr_lg_div_88_62_n_87);
  gl_gr_lg_div_88_62_g3721 : AOI21D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_80, A2 => gl_gr_lg_div_88_62_n_55, B => gl_gr_lg_div_88_62_n_75, ZN => gl_gr_lg_div_88_62_n_86);
  gl_gr_lg_div_88_62_g3722 : MAOI22D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_77, A2 => gl_n_92, B1 => gl_gr_lg_div_88_62_n_77, B2 => gl_n_92, ZN => gl_gr_lg_div_88_62_n_85);
  gl_gr_lg_div_88_62_g3723 : IND2D1BWP7T port map(A1 => gl_gr_lg_div_88_62_n_77, B1 => gl_n_92, ZN => gl_gr_lg_div_88_62_n_84);
  gl_gr_lg_div_88_62_g3724 : AOI21D0BWP7T port map(A1 => gl_n_92, A2 => gl_n_91, B => gl_gr_lg_div_88_62_n_76, ZN => gl_gr_lg_div_88_62_n_83);
  gl_gr_lg_div_88_62_g3725 : INVD0BWP7T port map(I => gl_gr_lg_div_88_62_n_82, ZN => gl_gr_lg_div_88_62_n_81);
  gl_gr_lg_div_88_62_g3726 : AOI221D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_70, A2 => gl_gr_lg_div_88_62_n_2, B1 => gl_gr_lg_div_88_62_n_66, B2 => gl_gr_lg_div_88_62_n_15, C => gl_gr_lg_div_88_62_n_73, ZN => gl_gr_lg_div_88_62_n_82);
  gl_gr_lg_div_88_62_g3727 : AO221D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_70, A2 => gl_gr_lg_div_88_62_n_63, B1 => gl_gr_lg_div_88_62_n_66, B2 => gl_gr_lg_div_88_62_n_59, C => gl_gr_lg_div_88_62_n_64, Z => gl_gr_lg_div_88_62_n_80);
  gl_gr_lg_div_88_62_g3728 : INVD0BWP7T port map(I => gl_gr_lg_div_88_62_n_78, ZN => gl_gr_lg_div_88_62_n_79);
  gl_gr_lg_div_88_62_g3729 : AOI221D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_70, A2 => gl_gr_lg_div_88_62_n_62, B1 => gl_gr_lg_div_88_62_n_64, B2 => gl_gr_lg_div_88_62_n_52, C => gl_gr_lg_div_88_62_n_74, ZN => gl_gr_lg_div_88_62_n_78);
  gl_gr_lg_div_88_62_g3730 : INVD0BWP7T port map(I => gl_gr_lg_div_88_62_n_77, ZN => gl_gr_lg_div_88_62_n_76);
  gl_gr_lg_div_88_62_g3731 : MAOI22D0BWP7T port map(A1 => gl_n_88, A2 => gl_gr_lg_div_88_62_n_7, B1 => gl_n_88, B2 => gl_gr_lg_div_88_62_n_7, ZN => gl_gr_lg_div_88_62_n_77);
  gl_gr_lg_div_88_62_g3732 : OAI32D1BWP7T port map(A1 => gl_gr_lg_div_88_62_n_55, A2 => gl_gr_lg_div_88_62_n_57, A3 => gl_gr_lg_div_88_62_n_71, B1 => gl_gr_lg_div_88_62_n_65, B2 => gl_gr_lg_div_88_62_n_69, ZN => gl_gr_lg_div_88_62_n_75);
  gl_gr_lg_div_88_62_g3733 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_71, A2 => gl_gr_lg_div_88_62_n_67, B1 => gl_gr_lg_div_88_62_n_66, B2 => gl_gr_lg_div_88_62_n_60, ZN => gl_gr_lg_div_88_62_n_74);
  gl_gr_lg_div_88_62_g3734 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_71, A2 => gl_gr_lg_div_88_62_n_15, B1 => gl_gr_lg_div_88_62_n_64, B2 => gl_n_94, ZN => gl_gr_lg_div_88_62_n_73);
  gl_gr_lg_div_88_62_g3735 : IND2D1BWP7T port map(A1 => gl_gr_lg_div_88_62_n_66, B1 => gl_gr_lg_div_88_62_n_71, ZN => gl_n_88);
  gl_gr_lg_div_88_62_g3736 : IND2D1BWP7T port map(A1 => gl_gr_lg_div_88_62_n_64, B1 => gl_gr_lg_div_88_62_n_68, ZN => gl_gr_lg_div_88_62_n_71);
  gl_gr_lg_div_88_62_g3737 : INVD0BWP7T port map(I => gl_gr_lg_div_88_62_n_70, ZN => gl_gr_lg_div_88_62_n_69);
  gl_gr_lg_div_88_62_g3738 : NR2D1BWP7T port map(A1 => gl_gr_lg_div_88_62_n_68, A2 => gl_gr_lg_div_88_62_n_66, ZN => gl_gr_lg_div_88_62_n_70);
  gl_gr_lg_div_88_62_g3739 : AOI21D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_65, A2 => gl_gr_lg_div_88_62_n_58, B => gl_gr_lg_div_88_62_n_61, ZN => gl_gr_lg_div_88_62_n_68);
  gl_gr_lg_div_88_62_g3740 : AOI21D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_63, A2 => gl_n_93, B => gl_gr_lg_div_88_62_n_57, ZN => gl_gr_lg_div_88_62_n_67);
  gl_gr_lg_div_88_62_g3741 : OA21D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_59, A2 => gl_gr_lg_div_88_62_n_55, B => gl_gr_lg_div_88_62_n_61, Z => gl_gr_lg_div_88_62_n_66);
  gl_gr_lg_div_88_62_g3742 : OR2D1BWP7T port map(A1 => gl_gr_lg_div_88_62_n_63, A2 => gl_gr_lg_div_88_62_n_55, Z => gl_gr_lg_div_88_62_n_65);
  gl_gr_lg_div_88_62_g3743 : AOI211XD0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_56, A2 => gl_gr_lg_div_88_62_n_55, B => gl_gr_lg_div_88_62_n_61, C => gl_gr_lg_div_88_62_n_58, ZN => gl_gr_lg_div_88_62_n_64);
  gl_gr_lg_div_88_62_g3744 : HA1D0BWP7T port map(A => gl_n_94, B => gl_gr_lg_div_88_62_n_52, CO => gl_gr_lg_div_88_62_n_63, S => gl_gr_lg_div_88_62_n_62);
  gl_gr_lg_div_88_62_g3745 : AO21D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_54, A2 => gl_gr_lg_div_88_62_n_31, B => gl_gr_lg_div_88_62_n_50, Z => gl_gr_lg_div_88_62_n_61);
  gl_gr_lg_div_88_62_g3746 : OAI21D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_51, A2 => gl_gr_lg_div_88_62_n_10, B => gl_gr_lg_div_88_62_n_59, ZN => gl_gr_lg_div_88_62_n_60);
  gl_gr_lg_div_88_62_g3747 : ND2D1BWP7T port map(A1 => gl_gr_lg_div_88_62_n_51, A2 => gl_gr_lg_div_88_62_n_10, ZN => gl_gr_lg_div_88_62_n_59);
  gl_gr_lg_div_88_62_g3748 : OAI21D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_47, A2 => gl_gr_lg_div_88_62_n_43, B => gl_gr_lg_div_88_62_n_53, ZN => gl_gr_lg_div_88_62_n_58);
  gl_gr_lg_div_88_62_g3749 : INVD0BWP7T port map(I => gl_gr_lg_div_88_62_n_56, ZN => gl_gr_lg_div_88_62_n_57);
  gl_gr_lg_div_88_62_g3750 : OAI21D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_2, A2 => gl_gr_lg_div_88_62_n_7, B => gl_gr_lg_div_88_62_n_51, ZN => gl_gr_lg_div_88_62_n_56);
  gl_gr_lg_div_88_62_g3751 : OAI221D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_45, A2 => gl_n_96, B1 => gl_gr_lg_div_88_62_n_14, B2 => gl_gr_lg_div_88_62_n_42, C => gl_gr_lg_div_88_62_n_49, ZN => gl_gr_lg_div_88_62_n_55);
  gl_gr_lg_div_88_62_g3752 : OAI221D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_45, A2 => gl_gr_lg_div_88_62_n_35, B1 => gl_gr_lg_div_88_62_n_39, B2 => gl_gr_lg_div_88_62_n_42, C => gl_gr_lg_div_88_62_n_40, ZN => gl_gr_lg_div_88_62_n_54);
  gl_gr_lg_div_88_62_g3753 : OA222D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_45, A2 => gl_gr_lg_div_88_62_n_37, B1 => gl_gr_lg_div_88_62_n_29, B2 => gl_gr_lg_div_88_62_n_40, C1 => gl_gr_lg_div_88_62_n_38, C2 => gl_gr_lg_div_88_62_n_42, Z => gl_gr_lg_div_88_62_n_53);
  gl_gr_lg_div_88_62_g3754 : INVD0BWP7T port map(I => gl_gr_lg_div_88_62_n_52, ZN => gl_gr_lg_div_88_62_n_51);
  gl_gr_lg_div_88_62_g3755 : MOAI22D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_48, A2 => gl_n_95, B1 => gl_gr_lg_div_88_62_n_48, B2 => gl_n_95, ZN => gl_gr_lg_div_88_62_n_52);
  gl_gr_lg_div_88_62_g3756 : OAI32D1BWP7T port map(A1 => gl_gr_lg_div_88_62_n_31, A2 => gl_gr_lg_div_88_62_n_34, A3 => gl_gr_lg_div_88_62_n_47, B1 => gl_gr_lg_div_88_62_n_41, B2 => gl_gr_lg_div_88_62_n_45, ZN => gl_gr_lg_div_88_62_n_50);
  gl_gr_lg_div_88_62_g3757 : MAOI22D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_46, A2 => gl_gr_lg_div_88_62_n_14, B1 => gl_gr_lg_div_88_62_n_40, B2 => gl_gr_lg_div_88_62_n_1, ZN => gl_gr_lg_div_88_62_n_49);
  gl_gr_lg_div_88_62_g3758 : INR2D1BWP7T port map(A1 => gl_gr_lg_div_88_62_n_42, B1 => gl_gr_lg_div_88_62_n_46, ZN => gl_gr_lg_div_88_62_n_48);
  gl_gr_lg_div_88_62_g3759 : INVD1BWP7T port map(I => gl_gr_lg_div_88_62_n_47, ZN => gl_gr_lg_div_88_62_n_46);
  gl_gr_lg_div_88_62_g3760 : ND2D1BWP7T port map(A1 => gl_gr_lg_div_88_62_n_44, A2 => gl_gr_lg_div_88_62_n_40, ZN => gl_gr_lg_div_88_62_n_47);
  gl_gr_lg_div_88_62_g3761 : IND2D1BWP7T port map(A1 => gl_gr_lg_div_88_62_n_44, B1 => gl_gr_lg_div_88_62_n_42, ZN => gl_gr_lg_div_88_62_n_45);
  gl_gr_lg_div_88_62_g3762 : AOI21D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_41, A2 => gl_gr_lg_div_88_62_n_32, B => gl_gr_lg_div_88_62_n_30, ZN => gl_gr_lg_div_88_62_n_44);
  gl_gr_lg_div_88_62_g3763 : IAO21D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_35, A2 => gl_gr_lg_div_88_62_n_3, B => gl_gr_lg_div_88_62_n_34, ZN => gl_gr_lg_div_88_62_n_43);
  gl_gr_lg_div_88_62_g3764 : OAI21D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_36, A2 => gl_gr_lg_div_88_62_n_31, B => gl_gr_lg_div_88_62_n_30, ZN => gl_gr_lg_div_88_62_n_42);
  gl_gr_lg_div_88_62_g3765 : IND2D1BWP7T port map(A1 => gl_gr_lg_div_88_62_n_31, B1 => gl_gr_lg_div_88_62_n_35, ZN => gl_gr_lg_div_88_62_n_41);
  gl_gr_lg_div_88_62_g3766 : AO211D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_33, A2 => gl_gr_lg_div_88_62_n_31, B => gl_gr_lg_div_88_62_n_32, C => gl_gr_lg_div_88_62_n_30, Z => gl_gr_lg_div_88_62_n_40);
  gl_gr_lg_div_88_62_g3767 : INVD0BWP7T port map(I => gl_gr_lg_div_88_62_n_36, ZN => gl_gr_lg_div_88_62_n_39);
  gl_gr_lg_div_88_62_g3768 : OA21D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_29, A2 => gl_gr_lg_div_88_62_n_11, B => gl_gr_lg_div_88_62_n_36, Z => gl_gr_lg_div_88_62_n_38);
  gl_gr_lg_div_88_62_g3769 : MAOI22D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_29, A2 => gl_n_96, B1 => gl_gr_lg_div_88_62_n_29, B2 => gl_n_96, ZN => gl_gr_lg_div_88_62_n_37);
  gl_gr_lg_div_88_62_g3770 : ND2D1BWP7T port map(A1 => gl_gr_lg_div_88_62_n_29, A2 => gl_gr_lg_div_88_62_n_11, ZN => gl_gr_lg_div_88_62_n_36);
  gl_gr_lg_div_88_62_g3771 : OR2D1BWP7T port map(A1 => gl_gr_lg_div_88_62_n_29, A2 => gl_gr_lg_div_88_62_n_1, Z => gl_gr_lg_div_88_62_n_35);
  gl_gr_lg_div_88_62_g3772 : INVD0BWP7T port map(I => gl_gr_lg_div_88_62_n_33, ZN => gl_gr_lg_div_88_62_n_34);
  gl_gr_lg_div_88_62_g3773 : OAI21D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_1, A2 => gl_gr_lg_div_88_62_n_3, B => gl_gr_lg_div_88_62_n_29, ZN => gl_gr_lg_div_88_62_n_33);
  gl_gr_lg_div_88_62_g3774 : OAI222D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_27, A2 => gl_gr_lg_div_88_62_n_23, B1 => gl_gr_lg_div_88_62_n_8, B2 => gl_gr_lg_div_88_62_n_25, C1 => gl_gr_lg_div_88_62_n_19, C2 => gl_gr_lg_div_88_62_n_24, ZN => gl_gr_lg_div_88_62_n_32);
  gl_gr_lg_div_88_62_g3775 : OAI222D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_27, A2 => gl_gr_lg_div_88_62_n_18, B1 => gl_gr_lg_div_88_62_n_6, B2 => gl_gr_lg_div_88_62_n_25, C1 => gl_n_98, C2 => gl_gr_lg_div_88_62_n_24, ZN => gl_gr_lg_div_88_62_n_31);
  gl_gr_lg_div_88_62_g3776 : OAI31D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_22, A2 => gl_n_100, A3 => gl_gr_lg_div_88_62_n_27, B => gl_gr_lg_div_88_62_n_28, ZN => gl_gr_lg_div_88_62_n_30);
  gl_gr_lg_div_88_62_g3777 : MAOI22D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_27, A2 => gl_n_97, B1 => gl_gr_lg_div_88_62_n_27, B2 => gl_n_97, ZN => gl_gr_lg_div_88_62_n_29);
  gl_gr_lg_div_88_62_g3778 : ND2D1BWP7T port map(A1 => gl_gr_lg_div_88_62_n_26, A2 => gl_n_100, ZN => gl_gr_lg_div_88_62_n_28);
  gl_gr_lg_div_88_62_g3779 : ND2D1BWP7T port map(A1 => gl_gr_lg_div_88_62_n_24, A2 => gl_gr_lg_div_88_62_n_25, ZN => gl_gr_lg_div_88_62_n_27);
  gl_gr_lg_div_88_62_g3780 : OAI21D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_24, A2 => gl_gr_lg_div_88_62_n_20, B => gl_gr_lg_div_88_62_n_25, ZN => gl_gr_lg_div_88_62_n_26);
  gl_gr_lg_div_88_62_g3781 : AO21D0BWP7T port map(A1 => gl_n_100, A2 => gl_gr_lg_div_88_62_n_21, B => gl_n_101, Z => gl_gr_lg_div_88_62_n_25);
  gl_gr_lg_div_88_62_g3782 : OAI21D0BWP7T port map(A1 => gl_n_100, A2 => gl_gr_lg_div_88_62_n_9, B => gl_n_101, ZN => gl_gr_lg_div_88_62_n_24);
  gl_gr_lg_div_88_62_g3783 : AOI21D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_9, A2 => gl_n_97, B => gl_gr_lg_div_88_62_n_22, ZN => gl_gr_lg_div_88_62_n_23);
  gl_gr_lg_div_88_62_g3784 : INVD1BWP7T port map(I => gl_gr_lg_div_88_62_n_22, ZN => gl_gr_lg_div_88_62_n_21);
  gl_gr_lg_div_88_62_g3785 : AOI21D0BWP7T port map(A1 => gl_n_98, A2 => gl_n_97, B => gl_n_99, ZN => gl_gr_lg_div_88_62_n_22);
  gl_gr_lg_div_88_62_g3786 : INVD0BWP7T port map(I => gl_gr_lg_div_88_62_n_9, ZN => gl_gr_lg_div_88_62_n_20);
  gl_gr_lg_div_88_62_g3787 : AOI22D0BWP7T port map(A1 => gl_n_99, A2 => gl_gr_lg_div_88_62_n_6, B1 => gl_gr_lg_div_88_62_n_8, B2 => gl_n_98, ZN => gl_gr_lg_div_88_62_n_19);
  gl_gr_lg_div_88_62_g3788 : MAOI22D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_6, A2 => gl_n_97, B1 => gl_gr_lg_div_88_62_n_6, B2 => gl_n_97, ZN => gl_gr_lg_div_88_62_n_18);
  gl_gr_lg_div_88_62_g3789 : MOAI22D0BWP7T port map(A1 => gl_n_90, A2 => gl_gr_lg_div_88_62_n_5, B1 => gl_n_90, B2 => gl_gr_lg_div_88_62_n_5, ZN => gl_gr_lg_div_88_62_n_17);
  gl_gr_lg_div_88_62_g3790 : MOAI22D0BWP7T port map(A1 => gl_n_92, A2 => gl_gr_lg_div_88_62_n_4, B1 => gl_n_92, B2 => gl_gr_lg_div_88_62_n_4, ZN => gl_gr_lg_div_88_62_n_16);
  gl_gr_lg_div_88_62_g3791 : AOI22D0BWP7T port map(A1 => gl_n_94, A2 => gl_gr_lg_div_88_62_n_7, B1 => gl_gr_lg_div_88_62_n_2, B2 => gl_n_93, ZN => gl_gr_lg_div_88_62_n_15);
  gl_gr_lg_div_88_62_g3792 : OAI22D0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_1, A2 => gl_n_95, B1 => gl_n_96, B2 => gl_gr_lg_div_88_62_n_3, ZN => gl_gr_lg_div_88_62_n_14);
  gl_gr_lg_div_88_62_g3793 : NR2D1BWP7T port map(A1 => gl_n_90, A2 => gl_n_89, ZN => gl_gr_lg_div_88_62_n_13);
  gl_gr_lg_div_88_62_g3794 : NR2D1BWP7T port map(A1 => gl_n_92, A2 => gl_n_91, ZN => gl_gr_lg_div_88_62_n_12);
  gl_gr_lg_div_88_62_g3795 : NR2XD0BWP7T port map(A1 => gl_n_96, A2 => gl_n_95, ZN => gl_gr_lg_div_88_62_n_11);
  gl_gr_lg_div_88_62_g3796 : NR2D1BWP7T port map(A1 => gl_n_94, A2 => gl_n_93, ZN => gl_gr_lg_div_88_62_n_10);
  gl_gr_lg_div_88_62_g3797 : NR2XD0BWP7T port map(A1 => gl_gr_lg_div_88_62_n_8, A2 => gl_gr_lg_div_88_62_n_6, ZN => gl_gr_lg_div_88_62_n_9);
  gl_gr_lg_div_88_62_g3798 : INVD0BWP7T port map(I => gl_n_99, ZN => gl_gr_lg_div_88_62_n_8);
  gl_gr_lg_div_88_62_g3799 : INVD1BWP7T port map(I => gl_n_93, ZN => gl_gr_lg_div_88_62_n_7);
  gl_gr_lg_div_88_62_g3800 : INVD1BWP7T port map(I => gl_n_98, ZN => gl_gr_lg_div_88_62_n_6);
  gl_gr_lg_div_88_62_g3801 : INVD1BWP7T port map(I => gl_n_89, ZN => gl_gr_lg_div_88_62_n_5);
  gl_gr_lg_div_88_62_g3802 : INVD1BWP7T port map(I => gl_n_91, ZN => gl_gr_lg_div_88_62_n_4);
  gl_gr_lg_div_88_62_g3803 : INVD0BWP7T port map(I => gl_n_95, ZN => gl_gr_lg_div_88_62_n_3);
  gl_gr_lg_div_88_62_g3804 : INVD0BWP7T port map(I => gl_n_94, ZN => gl_gr_lg_div_88_62_n_2);
  gl_gr_lg_div_88_62_g3805 : INVD1BWP7T port map(I => gl_n_96, ZN => gl_gr_lg_div_88_62_n_1);
  ml_ms_ed_reg2_reg : DFQD1BWP7T port map(CP => CTS_20, D => FE_PHN53_ml_ms_ed_reg1, Q => ml_ms_ed_reg2);
  ml_ms_ed_g224 : NR2XD0BWP7T port map(A1 => ml_ms_ed_n_9, A2 => ml_ms_ed_state(0), ZN => ml_ms_output_edgedet);
  ml_ms_ed_g399 : OAI32D1BWP7T port map(A1 => FE_OFN35_reset, A2 => FE_PHN610_ml_ms_ed_state_1, A3 => FE_PHN547_ml_ms_ed_n_5, B1 => ml_ms_ed_n_9, B2 => ml_ms_ed_n_6, ZN => ml_ms_ed_n_8);
  ml_ms_ed_g400 : INVD0BWP7T port map(I => ml_ms_ed_n_6, ZN => ml_ms_ed_n_7);
  ml_ms_ed_g401 : IND2D1BWP7T port map(A1 => FE_OFN35_reset, B1 => FE_PHN547_ml_ms_ed_n_5, ZN => ml_ms_ed_n_6);
  ml_ms_ed_g402 : OAI31D0BWP7T port map(A1 => FE_PHN61_ml_ms_count_debounce_9, A2 => ml_ms_count_debounce(8), A3 => ml_ms_ed_n_4, B => ml_ms_ed_state(0), ZN => ml_ms_ed_n_5);
  ml_ms_ed_g403 : OR4D1BWP7T port map(A1 => FE_PHN123_ml_ms_count_debounce_11, A2 => FE_PHN433_ml_ms_count_debounce_10, A3 => FE_PHN615_ml_ms_count_debounce_12, A4 => ml_ms_ed_n_3, Z => ml_ms_ed_n_4);
  ml_ms_ed_g404 : OA31D1BWP7T port map(A1 => ml_ms_count_debounce(3), A2 => FE_PHN69_ml_ms_count_debounce_5, A3 => ml_ms_count_debounce(4), B => ml_ms_ed_n_1, Z => ml_ms_ed_n_3);
  ml_ms_ed_g405 : AO211D0BWP7T port map(A1 => ml_ms_ed_n_0, A2 => FE_PHN636_ml_ms_ed_reg2, B => FE_PHN610_ml_ms_ed_state_1, C => ml_ms_ed_state(0), Z => ml_ms_ed_n_2);
  ml_ms_ed_g406 : AN2D0BWP7T port map(A1 => FE_PHN513_ml_ms_count_debounce_6, A2 => FE_PHN473_ml_ms_count_debounce_7, Z => ml_ms_ed_n_1);
  ml_ms_ed_state_reg_0 : DFKCND1BWP7T port map(CN => FE_PHN621_ml_ms_ed_n_2, CP => CTS_20, D => ml_ms_ed_n_7, Q => FE_PHN614_ml_ms_ed_state_0, QN => ml_ms_count_debounce_reset);
  ml_ms_ed_state_reg_1 : DFD1BWP7T port map(CP => CTS_20, D => FE_PHN622_ml_ms_ed_n_8, Q => ml_ms_ed_state(1), QN => ml_ms_ed_n_9);
  ml_ms_ed_reg1_reg : DFD1BWP7T port map(CP => CTS_20, D => FE_PHN83_clk15k_in, Q => ml_ms_ed_reg1, QN => ml_ms_ed_n_0);

end routed;
