configuration countdown_bar_behav_cfg of countdown_bar is
   for behav
      for all: edge_det_fall use configuration work.edge_det_fall_behav_cfg;
      end for;
   end for;
end countdown_bar_behav_cfg;
