configuration submod_hcount_behaviour_cfg of submod_hcount is
   for behaviour
   end for;
end submod_hcount_behaviour_cfg;
